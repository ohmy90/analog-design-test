* NGSPICE file created from tt_um_ohmy90_ringOscillator.ext - technology: sky130B

.subckt sky130_fd_sc_hs__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM a_1100_75# a_1107_347#
+ a_318_389# a_315_75# a_916_347# a_69_260# a_936_75# a_465_249# a_237_75# a_501_75#
+ a_509_347# a_217_368#
X0 a_465_249# B a_936_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=3584,184
X1 a_501_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=6763,255 d=3584,184
X2 a_318_389# B a_217_368# VPB sky130_fd_pr__pfet_01v8 ad=0.19588 pd=1.565 as=0.18669 ps=1.46 w=1 l=0.15
**devattr s=7467,292 d=7835,313
X3 VPWR CIN a_509_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.1725 ps=1.345 w=1 l=0.15
**devattr s=7100,271 d=6200,262
X4 a_69_260# CIN a_315_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=4992,206
X5 a_501_75# a_465_249# a_69_260# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.1248 ps=1.03 w=0.64 l=0.15
**devattr s=4992,206 d=4608,200
X6 VGND A a_1100_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.29627 ps=1.75667 w=0.64 l=0.15
**devattr s=14384,346 d=8491,282
X7 VGND a_69_260# SUM VNB sky130_fd_pr__nfet_01v8_lvt ad=0.20595 pd=1.54456 as=0.2109 ps=2.05 w=0.74 l=0.15
**devattr s=8436,410 d=7663,279
X8 VGND CIN a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.1024 ps=0.96 w=0.64 l=0.15
**devattr s=3584,184 d=6336,227
X9 a_237_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=7663,279 d=3072,176
X10 a_509_347# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=9745,328 d=7100,271
X11 COUT a_465_249# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.26955 ps=1.84485 w=1.12 l=0.15
**devattr s=13216,566 d=12768,562
X12 a_465_249# B a_916_347# VPB sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1775 ps=1.355 w=1 l=0.15
**devattr s=7100,271 d=6000,260
X13 a_1107_347# CIN a_465_249# VPB sky130_fd_pr__pfet_01v8 ad=0.26 pd=1.85333 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6000,260 d=8900,289
X14 VPWR A a_1107_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.26 ps=1.85333 w=1 l=0.15
**devattr s=8900,289 d=13962,352
X15 COUT a_465_249# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.20595 ps=1.54456 w=0.74 l=0.15
**devattr s=7844,402 d=7992,404
X16 a_1100_75# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.29627 pd=1.75667 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=8491,282 d=6784,362
X17 a_509_347# a_465_249# a_69_260# VPB sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6000,260 d=6700,267
X18 a_217_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.18669 pd=1.46 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=7960,297 d=7467,292
X19 a_916_347# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1775 pd=1.355 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=6200,262 d=7100,271
X20 a_936_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=6336,227 d=3072,176
X21 a_69_260# CIN a_318_389# VPB sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.19588 ps=1.565 w=1 l=0.15
**devattr s=7835,313 d=6000,260
X22 a_1100_75# CIN a_465_249# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.29627 pd=1.75667 as=0.0896 ps=0.92 w=0.64 l=0.15
**devattr s=3584,184 d=14384,346
X23 VPWR a_69_260# SUM VPB sky130_fd_pr__pfet_01v8 ad=0.26955 pd=1.84485 as=0.3192 ps=2.81 w=1.12 l=0.15
**devattr s=12768,562 d=7960,297
X24 VPWR B a_509_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.1725 ps=1.345 w=1 l=0.15
**devattr s=6700,267 d=9745,328
X25 a_1107_347# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.26 pd=1.85333 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=13962,352 d=13400,534
X26 a_315_75# B a_237_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=3072,176
X27 VGND B a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.1024 ps=0.96 w=0.64 l=0.15
**devattr s=4608,200 d=6763,255
C0 a_1107_347# VPB 0.01475f
C1 VPB VPWR 0.24573f
C2 CIN B 0.19591f
C3 a_501_75# A 0.1337f
C4 a_1107_347# A 0.01477f
C5 VPB B 0.62725f
C6 VPWR A 0.04912f
C7 a_315_75# A 0.00252f
C8 VPWR a_509_347# 0.1543f
C9 B A 0.26846f
C10 SUM VPWR 0.10504f
C11 a_315_75# SUM 0
C12 VGND a_936_75# 0.0076f
C13 B a_509_347# 0.02783f
C14 B SUM 0
C15 CIN a_1100_75# 0.00368f
C16 a_69_260# a_936_75# 0
C17 A a_1100_75# 0.01955f
C18 a_237_75# VGND 0.00252f
C19 a_465_249# VGND 0.12651f
C20 COUT a_465_249# 0.06928f
C21 a_237_75# a_69_260# 0.00693f
C22 a_465_249# a_69_260# 0.03228f
C23 CIN a_318_389# 0.00717f
C24 a_501_75# VGND 0.14715f
C25 CIN VPB 0.12323f
C26 a_1107_347# VGND 0.00417f
C27 a_315_75# VGND 0.00207f
C28 VPWR VGND 0.08465f
C29 a_465_249# a_916_347# 0.0195f
C30 a_1107_347# COUT 0
C31 A a_217_368# 0
C32 CIN A 0.46738f
C33 COUT VPWR 0.12179f
C34 B VGND 0.04033f
C35 VPB A 0.14325f
C36 CIN a_509_347# 0.02394f
C37 COUT B 0.00688f
C38 CIN SUM 0
C39 a_501_75# a_69_260# 0.02578f
C40 VPWR a_69_260# 0.1278f
C41 a_315_75# a_69_260# 0.00702f
C42 VPB a_509_347# 0.00536f
C43 VPB SUM 0.01283f
C44 B a_69_260# 0.03966f
C45 A a_509_347# 0.01252f
C46 SUM A 0
C47 VGND a_1100_75# 0.25139f
C48 a_916_347# VPWR 0.01147f
C49 a_465_249# a_936_75# 0.00268f
C50 COUT a_1100_75# 0.00223f
C51 a_69_260# a_1100_75# 0
C52 a_237_75# a_465_249# 0
C53 a_501_75# a_936_75# 0
C54 VGND a_217_368# 0.0017f
C55 CIN VGND 0.13789f
C56 VPB VGND 0.01302f
C57 CIN COUT 0
C58 COUT VPB 0.01419f
C59 a_501_75# a_465_249# 0.00555f
C60 a_69_260# a_217_368# 0.01644f
C61 a_1107_347# a_465_249# 0.15034f
C62 A VGND 0.13151f
C63 a_237_75# VPWR 0
C64 a_315_75# a_465_249# 0
C65 a_465_249# VPWR 0.19408f
C66 CIN a_69_260# 0.10678f
C67 a_69_260# a_318_389# 0.02061f
C68 COUT A 0
C69 SUM VGND 0.0376f
C70 VPB a_69_260# 0.04981f
C71 B a_465_249# 0.27222f
C72 a_936_75# a_1100_75# 0
C73 A a_69_260# 0.27191f
C74 CIN a_916_347# 0.0061f
C75 a_69_260# a_509_347# 0.0624f
C76 SUM a_69_260# 0.12447f
C77 a_1107_347# VPWR 0.21905f
C78 a_916_347# A 0.0016f
C79 a_465_249# a_1100_75# 0.21113f
C80 a_501_75# B 0.00904f
C81 a_1107_347# B 0.06557f
C82 a_916_347# a_509_347# 0
C83 B VPWR 0.21956f
C84 CIN a_936_75# 0.00177f
C85 A a_936_75# 0.00492f
C86 VPWR a_1100_75# 0.00321f
C87 COUT VGND 0.07419f
C88 CIN a_465_249# 0.29824f
C89 B a_1100_75# 0.01175f
C90 a_465_249# a_318_389# 0
C91 VPB a_465_249# 0.10732f
C92 VGND a_69_260# 0.15999f
C93 a_237_75# A 0.00252f
C94 a_465_249# A 0.35643f
C95 a_465_249# a_509_347# 0.1366f
C96 a_237_75# SUM 0
C97 CIN a_501_75# 0.01116f
C98 VPWR a_217_368# 0.01541f
C99 a_1107_347# CIN 0.00192f
C100 CIN VPWR 0.13494f
C101 CIN a_315_75# 0.00121f
C102 VPWR a_318_389# 0.01234f
C103 VGND VNB 0.99802f
C104 COUT VNB 0.11284f
C105 CIN VNB 0.31573f
C106 A VNB 0.49885f
C107 VPWR VNB 0.79012f
C108 SUM VNB 0.11694f
C109 B VNB 0.61239f
C110 VPB VNB 2.08861f
C111 a_1100_75# VNB 0.01137f
C112 a_501_75# VNB 0.00504f
C113 a_1107_347# VNB 0.00204f
C114 a_509_347# VNB 0.00129f
C115 a_465_249# VNB 0.30402f
C116 a_69_260# VNB 0.15472f
.ends

.subckt sky130_fd_sc_hd__inv_6 a_37_47# w_n38_261# a_27_297# a_143_47# a_21_199# VSUBS
X0 a_27_297# a_21_199# a_143_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.20667 pd=1.74667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X1 a_143_47# a_21_199# a_27_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20667 ps=1.74667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 a_143_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12892 ps=1.26333 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X3 a_27_297# a_21_199# a_143_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.20667 pd=1.74667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 a_143_47# a_21_199# a_27_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20667 ps=1.74667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X5 a_27_297# a_21_199# a_143_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.20667 pd=1.74667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X6 a_143_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12892 ps=1.26333 w=0.65 l=0.15
**devattr s=9880,412 d=3510,184
X7 a_143_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12892 ps=1.26333 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X8 a_143_47# a_21_199# a_27_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20667 ps=1.74667 w=1 l=0.15
**devattr s=17200,572 d=5400,254
X9 a_37_47# a_21_199# a_143_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12892 pd=1.26333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X10 a_37_47# a_21_199# a_143_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12892 pd=1.26333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X11 a_37_47# a_21_199# a_143_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12892 pd=1.26333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=7020,368
C0 a_21_199# a_27_297# 0.13608f
C1 w_n38_261# a_21_199# 0.21261f
C2 a_37_47# a_21_199# 0.1215f
C3 a_143_47# a_27_297# 0.53032f
C4 a_143_47# w_n38_261# 0.01838f
C5 w_n38_261# a_27_297# 0.07832f
C6 a_143_47# a_37_47# 0.32587f
C7 a_37_47# a_27_297# 0.06953f
C8 a_37_47# w_n38_261# 0.00676f
C9 a_143_47# a_21_199# 0.54356f
C10 a_37_47# VSUBS 0.42142f
C11 a_143_47# VSUBS 0.09005f
C12 a_27_297# VSUBS 0.37325f
C13 a_21_199# VSUBS 0.64634f
C14 w_n38_261# VSUBS 0.69336f
.ends

.subckt sky130_fd_sc_hd__inv_4 a_37_47# w_n38_261# a_37_297# a_119_47# a_21_199# VSUBS
X0 a_37_297# a_21_199# a_119_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 a_119_47# a_21_199# a_37_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 a_119_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12837 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_37_297# a_21_199# a_119_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 a_37_47# a_21_199# a_119_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12837 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X5 a_119_47# a_21_199# a_37_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X6 a_37_47# a_21_199# a_119_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12837 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X7 a_119_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12837 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 a_21_199# a_37_297# 0.09823f
C1 w_n38_261# a_21_199# 0.14198f
C2 a_37_47# a_21_199# 0.08191f
C3 a_119_47# a_37_297# 0.36178f
C4 a_119_47# w_n38_261# 0.0159f
C5 w_n38_261# a_37_297# 0.06539f
C6 a_119_47# a_37_47# 0.26259f
C7 a_37_47# a_37_297# 0.05009f
C8 a_37_47# w_n38_261# 0.00667f
C9 a_119_47# a_21_199# 0.35989f
C10 a_37_47# VSUBS 0.32682f
C11 a_119_47# VSUBS 0.08495f
C12 a_37_297# VSUBS 0.29639f
C13 a_21_199# VSUBS 0.45186f
C14 w_n38_261# VSUBS 0.51617f
.ends

.subckt sky130_fd_sc_hd__inv_2 w_n38_261# a_111_47# a_29_47# a_21_199# a_29_297# VSUBS
X0 a_111_47# a_21_199# a_29_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1 a_29_47# a_21_199# a_111_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 a_111_47# a_21_199# a_29_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_29_297# a_21_199# a_111_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
C0 a_21_199# a_29_297# 0.06305f
C1 w_n38_261# a_21_199# 0.07418f
C2 a_29_47# a_21_199# 0.06375f
C3 a_111_47# a_29_297# 0.2091f
C4 a_111_47# w_n38_261# 0.0061f
C5 w_n38_261# a_29_297# 0.05206f
C6 a_111_47# a_29_47# 0.1546f
C7 a_29_47# a_29_297# 0.04227f
C8 a_29_47# w_n38_261# 0.00649f
C9 a_111_47# a_21_199# 0.08939f
C10 a_29_47# VSUBS 0.26619f
C11 a_111_47# VSUBS 0.03316f
C12 a_29_297# VSUBS 0.24604f
C13 a_21_199# VSUBS 0.26281f
C14 w_n38_261# VSUBS 0.33898f
.ends

.subckt sky130_fd_sc_hs__inv_2 a_114_368# w_n38_332# a_27_368# a_30_74# a_21_260#
+ VSUBS
X0 a_114_368# a_21_260# a_30_74# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
**devattr s=8436,410 d=4144,204
X1 a_27_368# a_21_260# a_114_368# w_n38_332# sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
**devattr s=6720,284 d=12768,562
X2 a_30_74# a_21_260# a_114_368# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
**devattr s=4144,204 d=8436,410
X3 a_114_368# a_21_260# a_27_368# w_n38_332# sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
**devattr s=12768,562 d=6720,284
C0 a_21_260# a_27_368# 0.07533f
C1 w_n38_332# a_21_260# 0.07759f
C2 a_30_74# a_21_260# 0.06173f
C3 a_114_368# a_27_368# 0.21165f
C4 a_114_368# w_n38_332# 0.00641f
C5 w_n38_332# a_27_368# 0.06315f
C6 a_114_368# a_30_74# 0.16424f
C7 a_30_74# a_27_368# 0.0376f
C8 a_30_74# w_n38_332# 0.00523f
C9 a_114_368# a_21_260# 0.11388f
C10 a_30_74# VSUBS 0.30324f
C11 a_114_368# VSUBS 0.04146f
C12 a_27_368# VSUBS 0.26758f
C13 a_21_260# VSUBS 0.30548f
C14 w_n38_332# VSUBS 0.40622f
.ends

.subckt sky130_fd_sc_hd__inv_1 a_150_47# w_n38_261# a_68_47# a_68_297# a_64_199# VSUBS
X0 a_150_47# a_64_199# a_68_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1 a_150_47# a_64_199# a_68_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
C0 a_64_199# a_68_297# 0.03703f
C1 w_n38_261# a_64_199# 0.04506f
C2 a_68_47# a_64_199# 0.04004f
C3 a_150_47# a_68_297# 0.12758f
C4 a_150_47# w_n38_261# 0.01774f
C5 w_n38_261# a_68_297# 0.05448f
C6 a_150_47# a_68_47# 0.09984f
C7 a_68_47# a_68_297# 0.03382f
C8 a_68_47# w_n38_261# 0.00948f
C9 a_150_47# a_64_199# 0.0476f
C10 a_68_47# VSUBS 0.25113f
C11 a_150_47# VSUBS 0.0961f
C12 a_68_297# VSUBS 0.21892f
C13 a_64_199# VSUBS 0.16664f
C14 w_n38_261# VSUBS 0.33898f
.ends

.subckt tt_um_ohmy90_ringOscillator clk A B CIN ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
Xsky130_fd_sc_hs__fa_1_6 A B sky130_fd_sc_hs__fa_1_6/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_4/CIN
+ SUM a_12918_2677# a_12925_2949# a_12136_2991# a_12133_2677# a_12734_2949# a_11902_3194#
+ a_12754_2677# a_13432_3194# a_12055_2677# a_12319_2677# a_12327_2949# a_12035_2970#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_7 A B sky130_fd_sc_hs__fa_1_7/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_6/CIN
+ SUM a_10856_2681# a_10863_2953# a_10074_2995# a_10071_2681# a_10672_2953# a_9840_3198#
+ a_10692_2681# a_11370_3198# a_9993_2681# a_10257_2681# a_10265_2953# a_9973_2974#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hd__inv_6_0 A sky130_fd_sc_hd__inv_6_0/w_n38_261# B ua[0] li_24174_2784#
+ VNB sky130_fd_sc_hd__inv_6
Xsky130_fd_sc_hd__inv_4_0 A sky130_fd_sc_hd__inv_4_0/w_n38_261# B li_24174_2784# li_23298_2790#
+ VNB sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/w_n38_261# li_23298_2790# A li_22720_2804#
+ B VNB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hs__fa_1_0 A B CIN A VNB VPB B sky130_fd_sc_hs__fa_1_1/CIN SUM a_2598_2695#
+ a_2605_2967# a_1816_3009# a_1813_2695# a_2414_2967# a_1582_3212# a_2434_2695# a_3112_3212#
+ a_1735_2695# a_1999_2695# a_2007_2967# a_1715_2988# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__inv_2_0 CIN sky130_fd_sc_hs__inv_2_0/w_n38_332# B A COUT VNB sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__fa_1_1 A B sky130_fd_sc_hs__fa_1_1/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_3/CIN
+ SUM a_4660_2691# a_4667_2963# a_3878_3005# a_3875_2691# a_4476_2963# a_3644_3208#
+ a_4496_2691# a_5174_3208# a_3797_2691# a_4061_2691# a_4069_2963# a_3777_2984# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hd__inv_1_0 li_22720_2804# sky130_fd_sc_hd__inv_1_0/w_n38_261# A B COUT
+ VNB sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hs__fa_1_2 A B sky130_fd_sc_hs__fa_1_2/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_7/CIN
+ SUM a_8796_2685# a_8803_2957# a_8014_2999# a_8011_2685# a_8612_2957# a_7780_3202#
+ a_8632_2685# a_9310_3202# a_7933_2685# a_8197_2685# a_8205_2957# a_7913_2978# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_4 A B sky130_fd_sc_hs__fa_1_4/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_5/CIN
+ SUM a_14992_2675# a_14999_2947# a_14210_2989# a_14207_2675# a_14808_2947# a_13976_3192#
+ a_14828_2675# a_15506_3192# a_14129_2675# a_14393_2675# a_14401_2947# a_14109_2968#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_3 A B sky130_fd_sc_hs__fa_1_3/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_2/CIN
+ SUM a_6734_2689# a_6741_2961# a_5952_3003# a_5949_2689# a_6550_2961# a_5718_3206#
+ a_6570_2689# a_7248_3206# a_5871_2689# a_6135_2689# a_6143_2961# a_5851_2982# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_5 A B sky130_fd_sc_hs__fa_1_5/CIN A VNB VPB B COUT SUM a_17054_2671#
+ a_17061_2943# a_16272_2985# a_16269_2671# a_16870_2943# a_16038_3188# a_16890_2671#
+ a_17568_3188# a_16191_2671# a_16455_2671# a_16463_2943# a_16171_2964# sky130_fd_sc_hs__fa_1
C0 a_13976_3192# a_14210_2989# -0
C1 a_5174_3208# a_3644_3208# 0
C2 a_4476_2963# A 0
C3 a_9840_3198# a_11370_3198# -0
C4 a_9840_3198# a_9310_3202# 0.00608f
C5 a_16455_2671# a_17568_3188# 0
C6 a_17568_3188# a_16870_2943# 0
C7 a_7780_3202# sky130_fd_sc_hs__fa_1_2/CIN 0.06636f
C8 B a_15506_3192# 0.04212f
C9 B sky130_fd_sc_hs__inv_2_0/w_n38_332# 0.01594f
C10 a_9310_3202# a_8612_2957# -0
C11 CIN A 0.20597f
C12 a_5174_3208# a_4496_2691# -0
C13 sky130_fd_sc_hs__fa_1_1/CIN a_3112_3212# 0.00578f
C14 a_11370_3198# sky130_fd_sc_hs__fa_1_7/CIN 0
C15 a_9310_3202# sky130_fd_sc_hs__fa_1_7/CIN 0.00636f
C16 li_24174_2784# A 0.11344f
C17 uio_out[6] uio_out[5] 0.03102f
C18 a_10265_2953# a_11370_3198# -0
C19 a_9310_3202# sky130_fd_sc_hs__fa_1_2/CIN 0
C20 a_7248_3206# A 0.02391f
C21 B a_8197_2685# 0.00184f
C22 VPB sky130_fd_sc_hs__fa_1_1/CIN 0.01675f
C23 sky130_fd_sc_hs__fa_1_1/CIN a_4667_2963# -0
C24 a_15506_3192# sky130_fd_sc_hs__fa_1_4/CIN 0
C25 sky130_fd_sc_hs__fa_1_5/CIN a_15506_3192# 0.00578f
C26 sky130_fd_sc_hs__fa_1_1/CIN a_4069_2963# 0
C27 B a_8014_2999# 0.00253f
C28 SUM a_9840_3198# 0
C29 B a_9973_2974# 0.00246f
C30 sky130_fd_sc_hd__inv_2_0/w_n38_261# COUT 0
C31 clk ena 0.03102f
C32 B a_12133_2677# 0
C33 a_13432_3194# COUT 0
C34 a_2598_2695# a_3112_3212# -0
C35 a_17054_2671# a_15506_3192# 0
C36 a_1813_2695# a_3112_3212# -0
C37 B a_12035_2970# 0.00246f
C38 a_7780_3202# A 0.00644f
C39 a_11370_3198# a_12918_2677# 0
C40 uio_out[6] uio_out[7] 0.03102f
C41 uo_out[4] uo_out[5] 0.03102f
C42 SUM sky130_fd_sc_hs__fa_1_7/CIN 0.07963f
C43 a_14401_2947# A 0.00225f
C44 a_7933_2685# sky130_fd_sc_hs__fa_1_2/CIN 0.00126f
C45 a_17568_3188# A 0.02392f
C46 B sky130_fd_sc_hd__inv_2_0/w_n38_261# 0.01331f
C47 a_4660_2691# CIN 0
C48 sky130_fd_sc_hs__fa_1_3/CIN a_5718_3206# 0.06234f
C49 B a_13432_3194# 0.04208f
C50 B a_14129_2675# -0
C51 a_13976_3192# COUT 0
C52 sky130_fd_sc_hs__fa_1_6/CIN a_12133_2677# 0
C53 SUM sky130_fd_sc_hs__fa_1_2/CIN 0.07889f
C54 sky130_fd_sc_hs__fa_1_6/CIN a_12035_2970# 0.00449f
C55 a_10257_2681# a_9840_3198# 0
C56 SUM sky130_fd_sc_hs__fa_1_3/CIN 0.07548f
C57 a_11370_3198# A 0.02406f
C58 a_9310_3202# A 0.02398f
C59 a_14207_2675# A 0
C60 a_16463_2943# A 0.00226f
C61 a_16269_2671# A 0
C62 B a_13976_3192# 0.00725f
C63 uio_oe[0] uio_out[7] 0.03102f
C64 a_3875_2691# A 0.00208f
C65 a_13432_3194# sky130_fd_sc_hs__fa_1_6/CIN 0
C66 a_10257_2681# sky130_fd_sc_hs__fa_1_7/CIN 0
C67 uo_out[0] uo_out[1] 0.03102f
C68 li_22720_2804# COUT 0.05798f
C69 B a_2007_2967# 0.0054f
C70 a_13432_3194# sky130_fd_sc_hs__fa_1_4/CIN 0.00595f
C71 sky130_fd_sc_hs__fa_1_4/CIN a_14129_2675# 0.00124f
C72 a_2414_2967# CIN 0.00304f
C73 a_5718_3206# A 0.00648f
C74 a_7933_2685# A 0
C75 B li_22720_2804# 0.08113f
C76 CIN COUT 0.07361f
C77 uio_out[4] uio_out[3] 0.03102f
C78 B a_14828_2675# 0
C79 a_5952_3003# CIN 0
C80 B a_3797_2691# -0
C81 B a_4476_2963# 0.00311f
C82 a_13976_3192# sky130_fd_sc_hs__fa_1_4/CIN 0.06234f
C83 a_5871_2689# CIN 0
C84 SUM A 0.02115f
C85 VPB a_15506_3192# 0
C86 li_24174_2784# COUT 0
C87 CIN a_6734_2689# 0
C88 B CIN 0.56347f
C89 a_12319_2677# A 0.0086f
C90 B li_24174_2784# 0.1041f
C91 a_13432_3194# a_11902_3194# 0
C92 a_14828_2675# sky130_fd_sc_hs__fa_1_4/CIN -0
C93 a_16038_3188# A 0.00658f
C94 a_7248_3206# a_6734_2689# -0
C95 B a_7248_3206# 0.04252f
C96 a_10257_2681# A 0.00859f
C97 a_12925_2949# A 0
C98 sky130_fd_sc_hs__fa_1_3/CIN a_6143_2961# 0
C99 a_3777_2984# sky130_fd_sc_hs__fa_1_1/CIN 0.00449f
C100 sky130_fd_sc_hs__fa_1_3/CIN a_6570_2689# -0
C101 a_17568_3188# COUT 0.02199f
C102 a_1816_3009# A 0.00186f
C103 uio_oe[5] uio_oe[4] 0.03102f
C104 B a_7780_3202# 0.00739f
C105 ua[0] sky130_fd_sc_hd__inv_4_0/w_n38_261# 0
C106 a_7913_2978# CIN 0
C107 a_12734_2949# A 0
C108 B a_14401_2947# 0.00607f
C109 a_11370_3198# COUT 0
C110 a_3644_3208# A 0.05965f
C111 a_9310_3202# COUT 0
C112 a_13432_3194# VPB 0
C113 B a_17568_3188# 0.04177f
C114 li_23298_2790# sky130_fd_sc_hd__inv_2_0/w_n38_261# 0.00671f
C115 sky130_fd_sc_hs__fa_1_1/CIN a_3878_3005# 0
C116 a_2007_2967# a_3112_3212# -0
C117 CIN a_6741_2961# 0.00105f
C118 sky130_fd_sc_hd__inv_1_0/w_n38_261# A 0.00166f
C119 a_4496_2691# A 0.00404f
C120 B a_11370_3198# 0.04232f
C121 B a_9310_3202# 0.04239f
C122 a_8632_2685# sky130_fd_sc_hs__fa_1_2/CIN -0
C123 sky130_fd_sc_hs__fa_1_3/CIN a_5851_2982# 0.0045f
C124 B a_14207_2675# 0
C125 a_6143_2961# A 0.00221f
C126 VPB a_13976_3192# 0
C127 B a_16463_2943# 0.00615f
C128 B a_16269_2671# 0
C129 ua[0] sky130_fd_sc_hd__inv_6_0/w_n38_261# 0.00885f
C130 B a_3875_2691# 0
C131 sky130_fd_sc_hs__fa_1_1/CIN a_2598_2695# -0
C132 uio_oe[2] uio_oe[3] 0.03102f
C133 a_6570_2689# A 0.00358f
C134 uo_out[6] uo_out[5] 0.03102f
C135 a_14401_2947# sky130_fd_sc_hs__fa_1_4/CIN 0
C136 uo_out[0] uio_in[7] 0.03102f
C137 sky130_fd_sc_hs__fa_1_5/CIN a_17568_3188# 0
C138 a_5871_2689# a_5718_3206# -0
C139 sky130_fd_sc_hs__fa_1_6/CIN a_11370_3198# 0.00642f
C140 CIN a_3112_3212# 0.03236f
C141 a_8205_2957# sky130_fd_sc_hs__fa_1_2/CIN 0
C142 a_8796_2685# sky130_fd_sc_hs__fa_1_7/CIN -0
C143 sky130_fd_sc_hs__fa_1_1/CIN a_2605_2967# 0
C144 B a_5718_3206# 0.00747f
C145 B a_7933_2685# -0
C146 a_10074_2995# sky130_fd_sc_hs__fa_1_7/CIN 0
C147 li_22720_2804# li_23298_2790# 0.05251f
C148 a_14207_2675# sky130_fd_sc_hs__fa_1_4/CIN 0
C149 a_4061_2691# a_5174_3208# 0
C150 sky130_fd_sc_hs__fa_1_5/CIN a_16463_2943# 0
C151 sky130_fd_sc_hs__fa_1_5/CIN a_16269_2671# 0
C152 a_8796_2685# sky130_fd_sc_hs__fa_1_2/CIN 0
C153 B SUM 0.02992f
C154 uio_out[3] uio_out[2] 0.03102f
C155 a_5851_2982# A -0
C156 a_1582_3212# a_1999_2695# 0
C157 a_2434_2695# CIN -0
C158 VPB CIN 0.03018f
C159 a_4667_2963# CIN 0.00106f
C160 a_8632_2685# A 0.00358f
C161 a_16038_3188# COUT 0
C162 a_5174_3208# sky130_fd_sc_hs__fa_1_3/CIN 0.00595f
C163 a_4069_2963# CIN 0.00118f
C164 B a_12319_2677# 0.00182f
C165 li_23298_2790# li_24174_2784# 0.03301f
C166 SUM sky130_fd_sc_hs__fa_1_6/CIN 0.07889f
C167 ua[0] A 0.03768f
C168 B a_16038_3188# 0.00716f
C169 VPB a_7248_3206# 0
C170 a_8205_2957# A 0.00222f
C171 B a_10257_2681# 0.00183f
C172 a_11370_3198# a_11902_3194# 0.00606f
C173 B a_12925_2949# 0.05134f
C174 a_14109_2968# A -0
C175 SUM sky130_fd_sc_hs__fa_1_4/CIN 0.07548f
C176 uo_out[6] uo_out[7] 0.03102f
C177 SUM sky130_fd_sc_hs__fa_1_5/CIN 0.07889f
C178 sky130_fd_sc_hs__fa_1_3/CIN a_6550_2961# 0
C179 sky130_fd_sc_hs__fa_1_6/CIN a_12319_2677# 0
C180 B a_1816_3009# 0.00221f
C181 a_8796_2685# A 0.01046f
C182 a_7780_3202# VPB 0
C183 a_10074_2995# A 0
C184 a_5174_3208# A 0.02785f
C185 B a_12734_2949# 0.0031f
C186 sky130_fd_sc_hs__fa_1_6/CIN a_12925_2949# -0
C187 sky130_fd_sc_hd__inv_1_0/w_n38_261# COUT 0.01108f
C188 VPB a_17568_3188# -0
C189 B a_3644_3208# 0.00746f
C190 sky130_fd_sc_hs__fa_1_5/CIN a_16038_3188# 0.06636f
C191 a_16890_2671# A 0.00359f
C192 sky130_fd_sc_hs__fa_1_4/CIN a_12925_2949# 0
C193 rst_n clk 0.03102f
C194 VPB a_11370_3198# 0.00733f
C195 B a_4496_2691# 0
C196 SUM a_11902_3194# 0
C197 B sky130_fd_sc_hd__inv_1_0/w_n38_261# 0.01507f
C198 VPB a_9310_3202# 0
C199 a_12734_2949# sky130_fd_sc_hs__fa_1_6/CIN 0
C200 B a_6143_2961# 0.00616f
C201 A a_6550_2961# 0
C202 a_14992_2675# A 0.01052f
C203 B a_6570_2689# 0
C204 SUM a_3112_3212# 0
C205 a_9840_3198# sky130_fd_sc_hs__fa_1_7/CIN 0.06628f
C206 uio_out[0] uo_out[7] 0.03102f
C207 a_1582_3212# A 0.01688f
C208 VPB a_5718_3206# 0
C209 a_5174_3208# a_4660_2691# -0
C210 sky130_fd_sc_hs__fa_1_2/CIN a_8612_2957# 0
C211 SUM VPB 0.01931f
C212 B a_5851_2982# 0.00243f
C213 uio_oe[6] uio_oe[7] 0.03102f
C214 a_12327_2949# a_13432_3194# 0
C215 sky130_fd_sc_hs__fa_1_7/CIN sky130_fd_sc_hs__fa_1_2/CIN -0
C216 a_3777_2984# CIN 0
C217 B a_8632_2685# 0
C218 a_10265_2953# sky130_fd_sc_hs__fa_1_7/CIN 0
C219 sky130_fd_sc_hs__fa_1_1/CIN a_3797_2691# 0.00126f
C220 uio_out[2] uio_out[1] 0.03102f
C221 sky130_fd_sc_hs__fa_1_1/CIN a_4476_2963# 0
C222 a_1999_2695# A 0.0099f
C223 sky130_fd_sc_hd__inv_4_0/w_n38_261# A 0.00128f
C224 VPB a_16038_3188# 0
C225 sky130_fd_sc_hs__fa_1_1/CIN CIN 0.00412f
C226 sky130_fd_sc_hs__fa_1_3/CIN sky130_fd_sc_hs__fa_1_2/CIN -0
C227 B ua[0] 0.03568f
C228 B a_8205_2957# 0.00624f
C229 a_14808_2947# A 0
C230 B a_14109_2968# 0.00241f
C231 a_3644_3208# a_3112_3212# 0.00606f
C232 a_8011_2685# sky130_fd_sc_hs__fa_1_2/CIN 0
C233 a_3878_3005# CIN 0
C234 a_9840_3198# A 0.0064f
C235 A a_8612_2957# 0
C236 a_16890_2671# COUT 0
C237 B a_8796_2685# 0.00714f
C238 ui_in[6] ui_in[7] 0.03102f
C239 a_5174_3208# a_6734_2689# 0
C240 ui_in[5] ui_in[4] 0.03102f
C241 B a_10074_2995# 0.00255f
C242 B a_5174_3208# 0.04248f
C243 sky130_fd_sc_hd__inv_6_0/w_n38_261# A 0
C244 sky130_fd_sc_hs__fa_1_7/CIN A 0.18163f
C245 a_14393_2675# A 0.00861f
C246 a_16870_2943# A 0
C247 a_16455_2671# A 0.00863f
C248 a_2598_2695# CIN 0
C249 VPB a_3644_3208# 0
C250 a_1735_2695# a_1582_3212# -0
C251 a_1715_2988# CIN 0.0017f
C252 a_4061_2691# A 0.07071f
C253 B a_16890_2671# 0
C254 a_14109_2968# sky130_fd_sc_hs__fa_1_4/CIN 0.0045f
C255 a_15506_3192# a_13976_3192# -0
C256 A sky130_fd_sc_hs__fa_1_2/CIN 0.17743f
C257 a_10265_2953# A 0.00223f
C258 sky130_fd_sc_hs__fa_1_3/CIN A 0.1782f
C259 a_10856_2681# a_11370_3198# -0
C260 a_2605_2967# CIN 0.00385f
C261 li_23298_2790# sky130_fd_sc_hd__inv_1_0/w_n38_261# 0
C262 a_10856_2681# a_9310_3202# 0
C263 a_10692_2681# sky130_fd_sc_hs__fa_1_7/CIN -0
C264 B a_6550_2961# 0.00307f
C265 a_8011_2685# A 0
C266 B a_14992_2675# 0.00709f
C267 A a_12918_2677# 0.0105f
C268 a_5949_2689# CIN 0
C269 sky130_fd_sc_hs__fa_1_7/CIN a_10863_2953# -0
C270 sky130_fd_sc_hs__fa_1_5/CIN a_16890_2671# -0
C271 a_6135_2689# CIN 0
C272 a_3875_2691# sky130_fd_sc_hs__fa_1_1/CIN 0
C273 B a_1582_3212# 0.01143f
C274 sky130_fd_sc_hs__inv_2_0/w_n38_332# CIN 0.0078f
C275 a_14992_2675# sky130_fd_sc_hs__fa_1_4/CIN 0
C276 a_6135_2689# a_7248_3206# 0
C277 sky130_fd_sc_hd__inv_4_0/w_n38_261# COUT 0
C278 sky130_fd_sc_hs__fa_1_3/CIN a_4660_2691# 0
C279 a_13432_3194# a_13976_3192# 0.00609f
C280 a_13976_3192# a_14129_2675# -0
C281 uio_oe[1] uio_oe[0] 0.03102f
C282 SUM sky130_fd_sc_hs__fa_1_1/CIN 0.07889f
C283 uio_in[2] uio_in[1] 0.03102f
C284 B a_1999_2695# 0.00187f
C285 a_9840_3198# COUT 0
C286 a_8197_2685# CIN 0
C287 a_10692_2681# A 0.00359f
C288 B sky130_fd_sc_hd__inv_4_0/w_n38_261# 0.0159f
C289 a_17061_2943# A 0
C290 ua[0] li_23298_2790# 0
C291 A a_14210_2989# 0
C292 uio_in[3] uio_in[2] 0.03102f
C293 a_8014_2999# CIN 0
C294 B a_14808_2947# 0.00306f
C295 li_22720_2804# sky130_fd_sc_hd__inv_2_0/w_n38_261# 0.00912f
C296 B a_9840_3198# 0.00738f
C297 a_10863_2953# A 0
C298 a_15506_3192# a_14401_2947# -0
C299 uio_in[4] uio_in[3] 0.03102f
C300 B a_8612_2957# 0.0031f
C301 a_4660_2691# A 0.01042f
C302 VPB a_5174_3208# 0
C303 B sky130_fd_sc_hs__fa_1_7/CIN 0.16279f
C304 B a_14393_2675# 0.00181f
C305 B sky130_fd_sc_hd__inv_6_0/w_n38_261# 0.00822f
C306 a_5174_3208# a_4069_2963# 0
C307 sky130_fd_sc_hs__fa_1_3/CIN a_5952_3003# 0
C308 B a_16870_2943# 0.00309f
C309 B a_16455_2671# 0.0018f
C310 B a_4061_2691# 0.00186f
C311 sky130_fd_sc_hd__inv_2_0/w_n38_261# li_24174_2784# 0
C312 sky130_fd_sc_hs__fa_1_3/CIN a_5871_2689# 0.00124f
C313 a_6734_2689# sky130_fd_sc_hs__fa_1_2/CIN -0
C314 a_14808_2947# sky130_fd_sc_hs__fa_1_4/CIN 0
C315 B sky130_fd_sc_hs__fa_1_2/CIN 0.16304f
C316 sky130_fd_sc_hs__fa_1_3/CIN a_6734_2689# 0
C317 B a_10265_2953# 0.00622f
C318 a_5949_2689# a_5718_3206# 0
C319 B sky130_fd_sc_hs__fa_1_3/CIN 0.17104f
C320 a_1735_2695# A 0.00107f
C321 sky130_fd_sc_hs__fa_1_6/CIN sky130_fd_sc_hs__fa_1_7/CIN -0
C322 sky130_fd_sc_hs__fa_1_1/CIN a_3644_3208# 0.06636f
C323 a_1582_3212# a_3112_3212# 0
C324 a_6135_2689# a_5718_3206# 0
C325 a_2007_2967# CIN 0.01499f
C326 B a_8011_2685# 0
C327 a_16171_2964# A -0
C328 a_14393_2675# sky130_fd_sc_hs__fa_1_4/CIN 0
C329 a_2414_2967# A 0.0014f
C330 sky130_fd_sc_hs__fa_1_5/CIN a_16870_2943# 0
C331 a_8197_2685# a_9310_3202# 0
C332 B a_12918_2677# 0.0071f
C333 sky130_fd_sc_hs__fa_1_5/CIN a_16455_2671# 0
C334 uio_oe[4] uio_oe[3] 0.03102f
C335 sky130_fd_sc_hs__fa_1_1/CIN a_4496_2691# -0
C336 A COUT 0.24319f
C337 a_5952_3003# A 0
C338 ui_in[0] rst_n 0.03102f
C339 VPB a_1582_3212# 0
C340 a_1582_3212# a_2434_2695# -0
C341 a_3797_2691# CIN 0
C342 SUM a_15506_3192# 0
C343 a_4476_2963# CIN 0
C344 a_5871_2689# A 0
C345 li_22720_2804# li_24174_2784# 0
C346 a_6734_2689# A 0.01043f
C347 sky130_fd_sc_hs__fa_1_6/CIN a_12918_2677# 0
C348 a_1999_2695# a_3112_3212# -0
C349 a_7913_2978# sky130_fd_sc_hs__fa_1_2/CIN 0.00449f
C350 B A 16.02574f
C351 uio_out[4] uio_out[5] 0.03102f
C352 a_12055_2677# A 0
C353 a_15506_3192# a_16038_3188# 0.00606f
C354 sky130_fd_sc_hs__fa_1_2/CIN a_6741_2961# 0
C355 sky130_fd_sc_hs__fa_1_3/CIN a_6741_2961# 0
C356 uio_in[7] uio_in[6] 0.03102f
C357 sky130_fd_sc_hs__fa_1_6/CIN A 0.1782f
C358 a_7248_3206# CIN 0.0035f
C359 a_12136_2991# A 0
C360 B a_10692_2681# 0
C361 sky130_fd_sc_hd__inv_4_0/w_n38_261# li_23298_2790# 0.00893f
C362 a_14207_2675# a_13976_3192# 0
C363 B a_17061_2943# 0.05131f
C364 B a_14210_2989# 0.00249f
C365 sky130_fd_sc_hs__fa_1_4/CIN A 0.17772f
C366 sky130_fd_sc_hs__fa_1_5/CIN A 0.1798f
C367 VPB a_9840_3198# 0
C368 a_7780_3202# CIN 0.00188f
C369 B a_10863_2953# 0.05137f
C370 a_17054_2671# A 0.01044f
C371 a_7913_2978# A -0
C372 SUM a_13432_3194# 0
C373 ui_in[0] ui_in[1] 0.03102f
C374 B a_4660_2691# 0.00717f
C375 VPB sky130_fd_sc_hs__fa_1_7/CIN 0.01694f
C376 sky130_fd_sc_hd__inv_6_0/w_n38_261# li_23298_2790# 0.00141f
C377 A a_6741_2961# 0
C378 a_17061_2943# sky130_fd_sc_hs__fa_1_5/CIN -0
C379 a_7780_3202# a_7248_3206# 0.00606f
C380 sky130_fd_sc_hs__fa_1_6/CIN a_10863_2953# 0
C381 SUM a_13976_3192# 0
C382 sky130_fd_sc_hs__fa_1_4/CIN a_14210_2989# 0
C383 a_13432_3194# a_12319_2677# 0
C384 VPB sky130_fd_sc_hs__fa_1_2/CIN 0.01668f
C385 a_9310_3202# CIN 0
C386 a_14999_2947# A 0
C387 a_5174_3208# sky130_fd_sc_hs__fa_1_1/CIN 0
C388 VPB sky130_fd_sc_hs__fa_1_3/CIN 0.01799f
C389 uio_in[1] uio_in[0] 0.03102f
C390 sky130_fd_sc_hs__fa_1_3/CIN a_4667_2963# 0
C391 B a_1735_2695# 0
C392 a_11902_3194# A 0.00651f
C393 a_3875_2691# CIN 0
C394 sky130_fd_sc_hs__fa_1_7/CIN a_8803_2957# 0
C395 a_12754_2677# A 0.00359f
C396 B a_16171_2964# 0.00245f
C397 B a_2414_2967# 0.00294f
C398 sky130_fd_sc_hs__fa_1_2/CIN a_8803_2957# -0
C399 a_3112_3212# A 0.02716f
C400 a_5718_3206# CIN 0.00192f
C401 a_7933_2685# CIN 0
C402 a_16272_2985# A 0
C403 B COUT 1.06958f
C404 B a_5952_3003# 0.00251f
C405 a_12734_2949# a_13432_3194# 0
C406 a_10672_2953# sky130_fd_sc_hs__fa_1_7/CIN 0
C407 B a_5871_2689# -0
C408 SUM CIN 0.0047f
C409 a_7780_3202# a_9310_3202# 0
C410 ui_in[2] ui_in[1] 0.03102f
C411 a_2434_2695# A 0.00384f
C412 B a_6734_2689# 0.00716f
C413 VPB A 0.03818f
C414 a_4667_2963# A 0
C415 li_23298_2790# A 0.11343f
C416 a_4069_2963# A 0.0022f
C417 a_7248_3206# a_5718_3206# 0
C418 sky130_fd_sc_hs__fa_1_5/CIN a_16171_2964# 0.00449f
C419 a_17568_3188# a_16463_2943# -0
C420 a_16269_2671# a_17568_3188# 0
C421 B a_12055_2677# -0
C422 SUM a_7248_3206# 0
C423 sky130_fd_sc_hs__fa_1_5/CIN COUT 0
C424 A a_8803_2957# 0
C425 B sky130_fd_sc_hs__fa_1_6/CIN 0.16326f
C426 B a_12136_2991# 0.00252f
C427 a_17054_2671# COUT 0.00121f
C428 a_4660_2691# a_3112_3212# 0
C429 SUM a_7780_3202# 0
C430 B sky130_fd_sc_hs__fa_1_4/CIN 0.16965f
C431 B sky130_fd_sc_hs__fa_1_5/CIN 0.16166f
C432 a_12055_2677# sky130_fd_sc_hs__fa_1_6/CIN 0.00126f
C433 a_1813_2695# a_1582_3212# 0
C434 a_1816_3009# CIN 0.00257f
C435 B a_17054_2671# 0.00708f
C436 B a_7913_2978# 0.00247f
C437 sky130_fd_sc_hs__fa_1_6/CIN a_12136_2991# 0
C438 a_10672_2953# A 0
C439 li_22720_2804# sky130_fd_sc_hd__inv_1_0/w_n38_261# 0.00934f
C440 a_1735_2695# a_3112_3212# 0
C441 a_3644_3208# CIN 0.00209f
C442 uio_in[4] uio_in[5] 0.03102f
C443 sky130_fd_sc_hs__fa_1_6/CIN sky130_fd_sc_hs__fa_1_4/CIN -0
C444 SUM a_11370_3198# 0
C445 a_10856_2681# sky130_fd_sc_hs__fa_1_7/CIN 0
C446 a_11902_3194# COUT 0
C447 SUM a_9310_3202# 0
C448 B a_6741_2961# 0.05141f
C449 ui_in[3] ui_in[2] 0.03102f
C450 a_4496_2691# CIN 0
C451 sky130_fd_sc_hs__fa_1_5/CIN sky130_fd_sc_hs__fa_1_4/CIN -0
C452 B a_14999_2947# 0.05133f
C453 a_17568_3188# a_16038_3188# 0
C454 a_6143_2961# CIN 0.00118f
C455 a_14992_2675# a_15506_3192# -0
C456 sky130_fd_sc_hs__fa_1_7/CIN a_9993_2681# 0.00127f
C457 B a_11902_3194# 0.00724f
C458 a_6570_2689# CIN 0
C459 sky130_fd_sc_hs__fa_1_5/CIN a_17054_2671# 0
C460 a_10071_2681# a_9840_3198# 0
C461 a_4061_2691# sky130_fd_sc_hs__fa_1_1/CIN 0
C462 B a_12754_2677# 0
C463 SUM a_5718_3206# 0
C464 sky130_fd_sc_hs__fa_1_3/CIN sky130_fd_sc_hs__fa_1_1/CIN -0
C465 a_10257_2681# a_11370_3198# 0
C466 B a_3112_3212# 0.04141f
C467 a_6143_2961# a_7248_3206# -0
C468 a_10071_2681# sky130_fd_sc_hs__fa_1_7/CIN 0
C469 uio_oe[6] uio_oe[5] 0.03102f
C470 sky130_fd_sc_hs__fa_1_6/CIN a_11902_3194# 0.06636f
C471 VPB COUT 0.0184f
C472 a_13976_3192# a_14109_2968# -0
C473 a_6570_2689# a_7248_3206# 0
C474 B a_16272_2985# 0.00251f
C475 li_23298_2790# COUT 0
C476 sky130_fd_sc_hs__fa_1_4/CIN a_14999_2947# 0
C477 a_12754_2677# sky130_fd_sc_hs__fa_1_6/CIN -0
C478 sky130_fd_sc_hs__fa_1_5/CIN a_14999_2947# 0
C479 a_5851_2982# CIN 0
C480 B a_2434_2695# 0
C481 B VPB 0.39719f
C482 B a_4667_2963# 0.05142f
C483 a_3777_2984# A -0
C484 ua[0] li_22720_2804# 0
C485 B li_23298_2790# 0.09658f
C486 a_10856_2681# A 0.01048f
C487 B a_4069_2963# 0.00628f
C488 a_16191_2671# A 0
C489 uio_in[0] ui_in[7] 0.03102f
C490 SUM a_16038_3188# 0
C491 ui_in[4] ui_in[3] 0.03102f
C492 a_14992_2675# a_13432_3194# 0
C493 sky130_fd_sc_hs__fa_1_1/CIN A 0.1836f
C494 a_9993_2681# A 0
C495 sky130_fd_sc_hs__fa_1_5/CIN a_16272_2985# 0
C496 VPB sky130_fd_sc_hs__fa_1_6/CIN 0.01661f
C497 B a_8803_2957# 0.05139f
C498 a_8205_2957# CIN 0
C499 ua[0] li_24174_2784# 0.03186f
C500 a_3878_3005# A 0
C501 VPB sky130_fd_sc_hs__fa_1_4/CIN 0.01809f
C502 sky130_fd_sc_hs__fa_1_5/CIN VPB 0.02401f
C503 a_5174_3208# a_4476_2963# -0
C504 a_10071_2681# A 0
C505 sky130_fd_sc_hs__fa_1_3/CIN a_5949_2689# 0
C506 a_14393_2675# a_15506_3192# 0
C507 SUM a_3644_3208# 0
C508 a_5174_3208# CIN 0.00351f
C509 uio_out[0] uio_out[1] 0.03102f
C510 sky130_fd_sc_hs__fa_1_3/CIN a_6135_2689# 0
C511 B a_10672_2953# 0.0031f
C512 a_2598_2695# A 0.01124f
C513 a_1715_2988# A 0.00175f
C514 a_1813_2695# A 0.00111f
C515 a_12327_2949# A 0.00224f
C516 uio_oe[2] uio_oe[1] 0.03102f
C517 a_8796_2685# a_7248_3206# 0
C518 a_9840_3198# a_9973_2974# 0
C519 a_2605_2967# A 0
C520 sky130_fd_sc_hs__fa_1_1/CIN a_4660_2691# 0
C521 VPB a_11902_3194# 0
C522 CIN a_6550_2961# 0
C523 sky130_fd_sc_hs__fa_1_7/CIN a_9973_2974# 0.00447f
C524 a_5949_2689# A 0
C525 a_8197_2685# sky130_fd_sc_hs__fa_1_2/CIN 0
C526 a_6135_2689# A 0.00856f
C527 a_2434_2695# a_3112_3212# 0
C528 VPB a_3112_3212# 0
C529 a_8014_2999# sky130_fd_sc_hs__fa_1_2/CIN 0
C530 a_1582_3212# CIN 0.00855f
C531 a_9310_3202# a_8205_2957# 0
C532 a_15506_3192# A 0.02417f
C533 sky130_fd_sc_hs__inv_2_0/w_n38_332# A 0
C534 a_8796_2685# a_9310_3202# -0
C535 a_16890_2671# a_17568_3188# -0
C536 li_22720_2804# sky130_fd_sc_hd__inv_4_0/w_n38_261# 0.00135f
C537 B a_3777_2984# 0.00247f
C538 B a_10856_2681# 0.00712f
C539 a_14393_2675# a_13976_3192# 0
C540 B a_16191_2671# -0
C541 uo_out[4] uo_out[3] 0.03102f
C542 a_1999_2695# CIN 0.00138f
C543 a_8197_2685# A 0.00857f
C544 B sky130_fd_sc_hs__fa_1_1/CIN 0.16275f
C545 B a_9993_2681# -0
C546 a_13432_3194# a_12918_2677# -0
C547 a_8014_2999# A 0
C548 a_5174_3208# a_5718_3206# 0.00609f
C549 a_10856_2681# sky130_fd_sc_hs__fa_1_6/CIN -0
C550 a_9973_2974# A -0
C551 A a_12133_2677# 0
C552 sky130_fd_sc_hd__inv_4_0/w_n38_261# li_24174_2784# 0.00648f
C553 li_22720_2804# sky130_fd_sc_hd__inv_6_0/w_n38_261# 0
C554 B a_3878_3005# 0.00253f
C555 a_12035_2970# A -0
C556 SUM a_5174_3208# 0
C557 uo_out[3] uo_out[2] 0.03102f
C558 B a_10071_2681# 0
C559 a_16191_2671# sky130_fd_sc_hs__fa_1_5/CIN 0.00126f
C560 sky130_fd_sc_hd__inv_2_0/w_n38_261# A 0.00177f
C561 a_13432_3194# A 0.02412f
C562 a_14129_2675# A 0
C563 B a_2598_2695# 0.00719f
C564 B a_1813_2695# 0
C565 B a_1715_2988# 0.00211f
C566 a_4061_2691# CIN 0
C567 sky130_fd_sc_hd__inv_6_0/w_n38_261# li_24174_2784# 0.01147f
C568 CIN sky130_fd_sc_hs__fa_1_2/CIN 0.00209f
C569 B a_12327_2949# 0.00619f
C570 uio_in[6] uio_in[5] 0.03102f
C571 a_13976_3192# A 0.00662f
C572 sky130_fd_sc_hs__fa_1_3/CIN CIN 0.00316f
C573 uo_out[2] uo_out[1] 0.03102f
C574 B a_2605_2967# 0.05145f
C575 a_2007_2967# A 0.0037f
C576 ui_in[6] ui_in[5] 0.03102f
C577 a_8011_2685# CIN 0
C578 a_7248_3206# sky130_fd_sc_hs__fa_1_2/CIN 0.00578f
C579 B a_5949_2689# 0
C580 a_12327_2949# sky130_fd_sc_hs__fa_1_6/CIN 0
C581 a_15506_3192# COUT 0
C582 SUM a_1582_3212# 0
C583 sky130_fd_sc_hs__fa_1_3/CIN a_7248_3206# 0
C584 sky130_fd_sc_hs__inv_2_0/w_n38_332# COUT 0.00689f
C585 li_22720_2804# A 0.08904f
C586 a_14828_2675# A 0.00359f
C587 B a_6135_2689# 0.00185f
C588 a_3797_2691# A 0.00202f
C589 ua[1] VNB 0.1369f
C590 ua[2] VNB 0.1369f
C591 ua[3] VNB 0.1369f
C592 ua[4] VNB 0.1369f
C593 ua[5] VNB 0.1369f
C594 ua[6] VNB 0.1369f
C595 ua[7] VNB 0.1369f
C596 ena VNB 0.06503f
C597 clk VNB 0.03887f
C598 rst_n VNB 0.03887f
C599 ui_in[0] VNB 0.03887f
C600 ui_in[1] VNB 0.03887f
C601 ui_in[2] VNB 0.03887f
C602 ui_in[3] VNB 0.03887f
C603 ui_in[4] VNB 0.03887f
C604 ui_in[5] VNB 0.03887f
C605 ui_in[6] VNB 0.03887f
C606 ui_in[7] VNB 0.03887f
C607 uio_in[0] VNB 0.03887f
C608 uio_in[1] VNB 0.03887f
C609 uio_in[2] VNB 0.03887f
C610 uio_in[3] VNB 0.03887f
C611 uio_in[4] VNB 0.03887f
C612 uio_in[5] VNB 0.03887f
C613 uio_in[6] VNB 0.03887f
C614 uio_in[7] VNB 0.03887f
C615 uo_out[0] VNB 0.03887f
C616 uo_out[1] VNB 0.03887f
C617 uo_out[2] VNB 0.03887f
C618 uo_out[3] VNB 0.03887f
C619 uo_out[4] VNB 0.03887f
C620 uo_out[5] VNB 0.03887f
C621 uo_out[6] VNB 0.03887f
C622 uo_out[7] VNB 0.03887f
C623 uio_out[0] VNB 0.03887f
C624 uio_out[1] VNB 0.03887f
C625 uio_out[2] VNB 0.03887f
C626 uio_out[3] VNB 0.03887f
C627 uio_out[4] VNB 0.03887f
C628 uio_out[5] VNB 0.03887f
C629 uio_out[6] VNB 0.03887f
C630 uio_out[7] VNB 0.03887f
C631 uio_oe[0] VNB 0.03887f
C632 uio_oe[1] VNB 0.03887f
C633 uio_oe[2] VNB 0.03887f
C634 uio_oe[3] VNB 0.03887f
C635 uio_oe[4] VNB 0.03887f
C636 uio_oe[5] VNB 0.03887f
C637 uio_oe[6] VNB 0.03887f
C638 uio_oe[7] VNB 0.06503f
C639 a_17568_3188# VNB 0.30402f
C640 a_16038_3188# VNB 0.14774f
C641 a_15506_3192# VNB 0.2969f
C642 a_13976_3192# VNB 0.14781f
C643 a_13432_3194# VNB 0.29703f
C644 a_11902_3194# VNB 0.14774f
C645 a_11370_3198# VNB 0.27898f
C646 a_9840_3198# VNB 0.1477f
C647 a_9310_3202# VNB 0.29686f
C648 a_7780_3202# VNB 0.14774f
C649 a_7248_3206# VNB 0.2969f
C650 a_5718_3206# VNB 0.14781f
C651 B VNB 27.75639f
C652 a_5174_3208# VNB 0.29703f
C653 a_3644_3208# VNB 0.14774f
C654 a_3112_3212# VNB 0.2969f
C655 CIN VNB 2.25303f
C656 a_1582_3212# VNB 0.15472f
C657 COUT VNB 4.95385f
C658 a_17054_2671# VNB 0.01137f
C659 a_16455_2671# VNB 0.00504f
C660 a_17061_2943# VNB 0.00204f
C661 a_16463_2943# VNB 0.00129f
C662 sky130_fd_sc_hs__fa_1_2/CIN VNB 0.44151f
C663 a_6734_2689# VNB 0.01137f
C664 a_6135_2689# VNB 0.00504f
C665 a_6741_2961# VNB 0.00204f
C666 a_6143_2961# VNB 0.00129f
C667 sky130_fd_sc_hs__fa_1_5/CIN VNB 0.32654f
C668 a_14992_2675# VNB 0.01137f
C669 a_14393_2675# VNB 0.00504f
C670 a_14999_2947# VNB 0.00204f
C671 a_14401_2947# VNB 0.00129f
C672 sky130_fd_sc_hs__fa_1_7/CIN VNB 0.44071f
C673 a_8796_2685# VNB 0.01137f
C674 a_8197_2685# VNB 0.00504f
C675 a_8803_2957# VNB 0.00204f
C676 a_8205_2957# VNB 0.00129f
C677 li_22720_2804# VNB 0.46538f
C678 sky130_fd_sc_hd__inv_1_0/w_n38_261# VNB 0.33898f
C679 sky130_fd_sc_hs__fa_1_3/CIN VNB 0.44533f
C680 a_4660_2691# VNB 0.01137f
C681 a_4061_2691# VNB 0.00504f
C682 a_4667_2963# VNB 0.00204f
C683 a_4069_2963# VNB 0.00129f
C684 sky130_fd_sc_hs__inv_2_0/w_n38_332# VNB 0.40622f
C685 sky130_fd_sc_hs__fa_1_1/CIN VNB 0.44129f
C686 A VNB 29.92727f
C687 SUM VNB 0.61793f
C688 VPB VNB 16.70885f
C689 a_2598_2695# VNB 0.01137f
C690 a_1999_2695# VNB 0.00504f
C691 a_2605_2967# VNB 0.00204f
C692 a_2007_2967# VNB 0.00129f
C693 sky130_fd_sc_hd__inv_2_0/w_n38_261# VNB 0.33898f
C694 li_24174_2784# VNB 0.84959f
C695 li_23298_2790# VNB 0.6013f
C696 sky130_fd_sc_hd__inv_4_0/w_n38_261# VNB 0.51617f
C697 ua[0] VNB 4.16862f
C698 sky130_fd_sc_hd__inv_6_0/w_n38_261# VNB 0.69336f
C699 sky130_fd_sc_hs__fa_1_6/CIN VNB 0.44099f
C700 a_10856_2681# VNB 0.01137f
C701 a_10257_2681# VNB 0.00504f
C702 a_10863_2953# VNB 0.00204f
C703 a_10265_2953# VNB 0.00129f
C704 sky130_fd_sc_hs__fa_1_4/CIN VNB 0.44615f
C705 a_12918_2677# VNB 0.01137f
C706 a_12319_2677# VNB 0.00504f
C707 a_12925_2949# VNB 0.00204f
C708 a_12327_2949# VNB 0.00129f
.ends

