magic
tech sky130B
magscale 1 2
timestamp 1752868562
<< nwell >>
rect 18084 5861 18436 6182
rect 26254 5813 27802 6134
rect 28060 5795 29608 6116
rect 1460 2952 3264 3324
rect 1798 2931 2994 2952
rect 3522 2948 5326 3320
rect 3860 2927 5056 2948
rect 5596 2946 7400 3318
rect 5934 2925 7130 2946
rect 7658 2942 9462 3314
rect 7996 2921 9192 2942
rect 9718 2938 11522 3310
rect 10056 2917 11252 2938
rect 11780 2934 13584 3306
rect 12118 2913 13314 2934
rect 13854 2932 15658 3304
rect 14192 2911 15388 2932
rect 15916 2928 17720 3300
rect 16254 2907 17450 2928
<< pwell >>
rect 18164 5621 18350 5803
rect 18164 5617 18185 5621
rect 18151 5583 18185 5617
rect 26306 5573 27752 5755
rect 26321 5535 26355 5573
rect 28112 5555 29558 5737
rect 28127 5517 28161 5555
rect 1499 2849 1688 2868
rect 3036 2849 3225 2868
rect 1499 2669 3225 2849
rect 3561 2845 3750 2864
rect 5098 2845 5287 2864
rect 1498 2620 3226 2669
rect 3561 2665 5287 2845
rect 5635 2843 5824 2862
rect 7172 2843 7361 2862
rect 3560 2616 5288 2665
rect 5635 2663 7361 2843
rect 7697 2839 7886 2858
rect 9234 2839 9423 2858
rect 5634 2614 7362 2663
rect 7697 2659 9423 2839
rect 9757 2835 9946 2854
rect 11294 2835 11483 2854
rect 7696 2610 9424 2659
rect 9757 2655 11483 2835
rect 11819 2831 12008 2850
rect 13356 2831 13545 2850
rect 9756 2606 11484 2655
rect 11819 2651 13545 2831
rect 13893 2829 14082 2848
rect 15430 2829 15619 2848
rect 11818 2602 13546 2651
rect 13893 2649 15619 2829
rect 15955 2825 16144 2844
rect 17492 2825 17681 2844
rect 13892 2600 15620 2649
rect 15955 2645 17681 2825
rect 15954 2596 17682 2645
<< nmoslvt >>
rect 1582 2694 1612 2842
rect 1705 2695 1735 2823
rect 1783 2695 1813 2823
rect 1861 2695 1891 2823
rect 1969 2695 1999 2823
rect 2071 2695 2101 2823
rect 2189 2695 2219 2823
rect 2275 2695 2305 2823
rect 2404 2695 2434 2823
rect 2482 2695 2512 2823
rect 2568 2695 2598 2823
rect 2780 2695 2810 2823
rect 2925 2695 2955 2823
rect 3115 2694 3145 2842
rect 3644 2690 3674 2838
rect 3767 2691 3797 2819
rect 3845 2691 3875 2819
rect 3923 2691 3953 2819
rect 4031 2691 4061 2819
rect 4133 2691 4163 2819
rect 4251 2691 4281 2819
rect 4337 2691 4367 2819
rect 4466 2691 4496 2819
rect 4544 2691 4574 2819
rect 4630 2691 4660 2819
rect 4842 2691 4872 2819
rect 4987 2691 5017 2819
rect 5177 2690 5207 2838
rect 5718 2688 5748 2836
rect 5841 2689 5871 2817
rect 5919 2689 5949 2817
rect 5997 2689 6027 2817
rect 6105 2689 6135 2817
rect 6207 2689 6237 2817
rect 6325 2689 6355 2817
rect 6411 2689 6441 2817
rect 6540 2689 6570 2817
rect 6618 2689 6648 2817
rect 6704 2689 6734 2817
rect 6916 2689 6946 2817
rect 7061 2689 7091 2817
rect 7251 2688 7281 2836
rect 7780 2684 7810 2832
rect 7903 2685 7933 2813
rect 7981 2685 8011 2813
rect 8059 2685 8089 2813
rect 8167 2685 8197 2813
rect 8269 2685 8299 2813
rect 8387 2685 8417 2813
rect 8473 2685 8503 2813
rect 8602 2685 8632 2813
rect 8680 2685 8710 2813
rect 8766 2685 8796 2813
rect 8978 2685 9008 2813
rect 9123 2685 9153 2813
rect 9313 2684 9343 2832
rect 9840 2680 9870 2828
rect 9963 2681 9993 2809
rect 10041 2681 10071 2809
rect 10119 2681 10149 2809
rect 10227 2681 10257 2809
rect 10329 2681 10359 2809
rect 10447 2681 10477 2809
rect 10533 2681 10563 2809
rect 10662 2681 10692 2809
rect 10740 2681 10770 2809
rect 10826 2681 10856 2809
rect 11038 2681 11068 2809
rect 11183 2681 11213 2809
rect 11373 2680 11403 2828
rect 11902 2676 11932 2824
rect 12025 2677 12055 2805
rect 12103 2677 12133 2805
rect 12181 2677 12211 2805
rect 12289 2677 12319 2805
rect 12391 2677 12421 2805
rect 12509 2677 12539 2805
rect 12595 2677 12625 2805
rect 12724 2677 12754 2805
rect 12802 2677 12832 2805
rect 12888 2677 12918 2805
rect 13100 2677 13130 2805
rect 13245 2677 13275 2805
rect 13435 2676 13465 2824
rect 13976 2674 14006 2822
rect 14099 2675 14129 2803
rect 14177 2675 14207 2803
rect 14255 2675 14285 2803
rect 14363 2675 14393 2803
rect 14465 2675 14495 2803
rect 14583 2675 14613 2803
rect 14669 2675 14699 2803
rect 14798 2675 14828 2803
rect 14876 2675 14906 2803
rect 14962 2675 14992 2803
rect 15174 2675 15204 2803
rect 15319 2675 15349 2803
rect 15509 2674 15539 2822
rect 16038 2670 16068 2818
rect 16161 2671 16191 2799
rect 16239 2671 16269 2799
rect 16317 2671 16347 2799
rect 16425 2671 16455 2799
rect 16527 2671 16557 2799
rect 16645 2671 16675 2799
rect 16731 2671 16761 2799
rect 16860 2671 16890 2799
rect 16938 2671 16968 2799
rect 17024 2671 17054 2799
rect 17236 2671 17266 2799
rect 17381 2671 17411 2799
rect 17571 2670 17601 2818
<< ndiff >>
rect 18190 5765 18242 5777
rect 18190 5731 18198 5765
rect 18232 5731 18242 5765
rect 18190 5697 18242 5731
rect 18190 5663 18198 5697
rect 18232 5663 18242 5697
rect 18190 5647 18242 5663
rect 18272 5765 18324 5777
rect 18272 5731 18282 5765
rect 18316 5731 18324 5765
rect 18272 5697 18324 5731
rect 18272 5663 18282 5697
rect 18316 5663 18324 5697
rect 18272 5647 18324 5663
rect 26332 5713 26384 5729
rect 26332 5679 26340 5713
rect 26374 5679 26384 5713
rect 26332 5645 26384 5679
rect 26332 5611 26340 5645
rect 26374 5611 26384 5645
rect 26332 5599 26384 5611
rect 26414 5713 26468 5729
rect 26414 5679 26424 5713
rect 26458 5679 26468 5713
rect 26414 5645 26468 5679
rect 26414 5611 26424 5645
rect 26458 5611 26468 5645
rect 26414 5599 26468 5611
rect 26498 5645 26552 5729
rect 26498 5611 26508 5645
rect 26542 5611 26552 5645
rect 26498 5599 26552 5611
rect 26582 5713 26636 5729
rect 26582 5679 26592 5713
rect 26626 5679 26636 5713
rect 26582 5645 26636 5679
rect 26582 5611 26592 5645
rect 26626 5611 26636 5645
rect 26582 5599 26636 5611
rect 26666 5645 26720 5729
rect 26666 5611 26676 5645
rect 26710 5611 26720 5645
rect 26666 5599 26720 5611
rect 26750 5713 26804 5729
rect 26750 5679 26760 5713
rect 26794 5679 26804 5713
rect 26750 5645 26804 5679
rect 26750 5611 26760 5645
rect 26794 5611 26804 5645
rect 26750 5599 26804 5611
rect 26834 5645 26888 5729
rect 26834 5611 26844 5645
rect 26878 5611 26888 5645
rect 26834 5599 26888 5611
rect 26918 5713 26972 5729
rect 26918 5679 26928 5713
rect 26962 5679 26972 5713
rect 26918 5645 26972 5679
rect 26918 5611 26928 5645
rect 26962 5611 26972 5645
rect 26918 5599 26972 5611
rect 27002 5645 27056 5729
rect 27002 5611 27012 5645
rect 27046 5611 27056 5645
rect 27002 5599 27056 5611
rect 27086 5713 27140 5729
rect 27086 5679 27096 5713
rect 27130 5679 27140 5713
rect 27086 5645 27140 5679
rect 27086 5611 27096 5645
rect 27130 5611 27140 5645
rect 27086 5599 27140 5611
rect 27170 5645 27224 5729
rect 27170 5611 27180 5645
rect 27214 5611 27224 5645
rect 27170 5599 27224 5611
rect 27254 5713 27308 5729
rect 27254 5679 27264 5713
rect 27298 5679 27308 5713
rect 27254 5645 27308 5679
rect 27254 5611 27264 5645
rect 27298 5611 27308 5645
rect 27254 5599 27308 5611
rect 27338 5645 27392 5729
rect 27338 5611 27348 5645
rect 27382 5611 27392 5645
rect 27338 5599 27392 5611
rect 27422 5713 27476 5729
rect 27422 5679 27432 5713
rect 27466 5679 27476 5713
rect 27422 5645 27476 5679
rect 27422 5611 27432 5645
rect 27466 5611 27476 5645
rect 27422 5599 27476 5611
rect 27506 5645 27560 5729
rect 27506 5611 27516 5645
rect 27550 5611 27560 5645
rect 27506 5599 27560 5611
rect 27590 5713 27644 5729
rect 27590 5679 27600 5713
rect 27634 5679 27644 5713
rect 27590 5645 27644 5679
rect 27590 5611 27600 5645
rect 27634 5611 27644 5645
rect 27590 5599 27644 5611
rect 27674 5713 27726 5729
rect 27674 5679 27684 5713
rect 27718 5679 27726 5713
rect 27674 5645 27726 5679
rect 27674 5611 27684 5645
rect 27718 5611 27726 5645
rect 27674 5599 27726 5611
rect 28138 5695 28190 5711
rect 28138 5661 28146 5695
rect 28180 5661 28190 5695
rect 28138 5627 28190 5661
rect 28138 5593 28146 5627
rect 28180 5593 28190 5627
rect 28138 5581 28190 5593
rect 28220 5695 28274 5711
rect 28220 5661 28230 5695
rect 28264 5661 28274 5695
rect 28220 5627 28274 5661
rect 28220 5593 28230 5627
rect 28264 5593 28274 5627
rect 28220 5581 28274 5593
rect 28304 5627 28358 5711
rect 28304 5593 28314 5627
rect 28348 5593 28358 5627
rect 28304 5581 28358 5593
rect 28388 5695 28442 5711
rect 28388 5661 28398 5695
rect 28432 5661 28442 5695
rect 28388 5627 28442 5661
rect 28388 5593 28398 5627
rect 28432 5593 28442 5627
rect 28388 5581 28442 5593
rect 28472 5627 28526 5711
rect 28472 5593 28482 5627
rect 28516 5593 28526 5627
rect 28472 5581 28526 5593
rect 28556 5695 28610 5711
rect 28556 5661 28566 5695
rect 28600 5661 28610 5695
rect 28556 5627 28610 5661
rect 28556 5593 28566 5627
rect 28600 5593 28610 5627
rect 28556 5581 28610 5593
rect 28640 5627 28694 5711
rect 28640 5593 28650 5627
rect 28684 5593 28694 5627
rect 28640 5581 28694 5593
rect 28724 5695 28778 5711
rect 28724 5661 28734 5695
rect 28768 5661 28778 5695
rect 28724 5627 28778 5661
rect 28724 5593 28734 5627
rect 28768 5593 28778 5627
rect 28724 5581 28778 5593
rect 28808 5627 28862 5711
rect 28808 5593 28818 5627
rect 28852 5593 28862 5627
rect 28808 5581 28862 5593
rect 28892 5695 28946 5711
rect 28892 5661 28902 5695
rect 28936 5661 28946 5695
rect 28892 5627 28946 5661
rect 28892 5593 28902 5627
rect 28936 5593 28946 5627
rect 28892 5581 28946 5593
rect 28976 5627 29030 5711
rect 28976 5593 28986 5627
rect 29020 5593 29030 5627
rect 28976 5581 29030 5593
rect 29060 5695 29114 5711
rect 29060 5661 29070 5695
rect 29104 5661 29114 5695
rect 29060 5627 29114 5661
rect 29060 5593 29070 5627
rect 29104 5593 29114 5627
rect 29060 5581 29114 5593
rect 29144 5627 29198 5711
rect 29144 5593 29154 5627
rect 29188 5593 29198 5627
rect 29144 5581 29198 5593
rect 29228 5695 29282 5711
rect 29228 5661 29238 5695
rect 29272 5661 29282 5695
rect 29228 5627 29282 5661
rect 29228 5593 29238 5627
rect 29272 5593 29282 5627
rect 29228 5581 29282 5593
rect 29312 5627 29366 5711
rect 29312 5593 29322 5627
rect 29356 5593 29366 5627
rect 29312 5581 29366 5593
rect 29396 5695 29450 5711
rect 29396 5661 29406 5695
rect 29440 5661 29450 5695
rect 29396 5627 29450 5661
rect 29396 5593 29406 5627
rect 29440 5593 29450 5627
rect 29396 5581 29450 5593
rect 29480 5695 29532 5711
rect 29480 5661 29490 5695
rect 29524 5661 29532 5695
rect 29480 5627 29532 5661
rect 29480 5593 29490 5627
rect 29524 5593 29532 5627
rect 29480 5581 29532 5593
rect 1525 2830 1582 2842
rect 1525 2796 1537 2830
rect 1571 2796 1582 2830
rect 1525 2740 1582 2796
rect 1525 2706 1537 2740
rect 1571 2706 1582 2740
rect 1525 2694 1582 2706
rect 1612 2823 1662 2842
rect 1612 2702 1705 2823
rect 1612 2694 1641 2702
rect 1627 2668 1641 2694
rect 1675 2695 1705 2702
rect 1735 2695 1783 2823
rect 1813 2695 1861 2823
rect 1891 2747 1969 2823
rect 1891 2713 1902 2747
rect 1936 2713 1969 2747
rect 1891 2695 1969 2713
rect 1999 2754 2071 2823
rect 1999 2720 2018 2754
rect 2052 2720 2071 2754
rect 1999 2695 2071 2720
rect 2101 2702 2189 2823
rect 2101 2695 2128 2702
rect 1675 2668 1690 2695
rect 1627 2656 1690 2668
rect 2116 2668 2128 2695
rect 2162 2695 2189 2702
rect 2219 2754 2275 2823
rect 2219 2720 2230 2754
rect 2264 2720 2275 2754
rect 2219 2695 2275 2720
rect 2305 2746 2404 2823
rect 2305 2712 2344 2746
rect 2378 2712 2404 2746
rect 2305 2695 2404 2712
rect 2434 2695 2482 2823
rect 2512 2757 2568 2823
rect 2512 2723 2523 2757
rect 2557 2723 2568 2757
rect 2512 2695 2568 2723
rect 2598 2705 2780 2823
rect 2598 2695 2625 2705
rect 2162 2668 2174 2695
rect 2613 2671 2625 2695
rect 2659 2671 2719 2705
rect 2753 2695 2780 2705
rect 2810 2698 2925 2823
rect 2810 2695 2864 2698
rect 2753 2671 2765 2695
rect 2116 2656 2174 2668
rect 2613 2659 2765 2671
rect 2852 2664 2864 2695
rect 2898 2695 2925 2698
rect 2955 2766 3008 2823
rect 2955 2732 2966 2766
rect 3000 2732 3008 2766
rect 2955 2695 3008 2732
rect 3062 2758 3115 2842
rect 3062 2724 3070 2758
rect 3104 2724 3115 2758
rect 2898 2664 2910 2695
rect 3062 2694 3115 2724
rect 3145 2830 3199 2842
rect 3145 2796 3156 2830
rect 3190 2796 3199 2830
rect 3145 2740 3199 2796
rect 3145 2706 3156 2740
rect 3190 2706 3199 2740
rect 3145 2694 3199 2706
rect 3587 2826 3644 2838
rect 3587 2792 3599 2826
rect 3633 2792 3644 2826
rect 3587 2736 3644 2792
rect 3587 2702 3599 2736
rect 3633 2702 3644 2736
rect 3587 2690 3644 2702
rect 3674 2819 3724 2838
rect 3674 2698 3767 2819
rect 3674 2690 3703 2698
rect 3689 2664 3703 2690
rect 3737 2691 3767 2698
rect 3797 2691 3845 2819
rect 3875 2691 3923 2819
rect 3953 2743 4031 2819
rect 3953 2709 3964 2743
rect 3998 2709 4031 2743
rect 3953 2691 4031 2709
rect 4061 2750 4133 2819
rect 4061 2716 4080 2750
rect 4114 2716 4133 2750
rect 4061 2691 4133 2716
rect 4163 2698 4251 2819
rect 4163 2691 4190 2698
rect 3737 2664 3752 2691
rect 2852 2656 2910 2664
rect 3689 2652 3752 2664
rect 4178 2664 4190 2691
rect 4224 2691 4251 2698
rect 4281 2750 4337 2819
rect 4281 2716 4292 2750
rect 4326 2716 4337 2750
rect 4281 2691 4337 2716
rect 4367 2742 4466 2819
rect 4367 2708 4406 2742
rect 4440 2708 4466 2742
rect 4367 2691 4466 2708
rect 4496 2691 4544 2819
rect 4574 2753 4630 2819
rect 4574 2719 4585 2753
rect 4619 2719 4630 2753
rect 4574 2691 4630 2719
rect 4660 2701 4842 2819
rect 4660 2691 4687 2701
rect 4224 2664 4236 2691
rect 4675 2667 4687 2691
rect 4721 2667 4781 2701
rect 4815 2691 4842 2701
rect 4872 2694 4987 2819
rect 4872 2691 4926 2694
rect 4815 2667 4827 2691
rect 4178 2652 4236 2664
rect 4675 2655 4827 2667
rect 4914 2660 4926 2691
rect 4960 2691 4987 2694
rect 5017 2762 5070 2819
rect 5017 2728 5028 2762
rect 5062 2728 5070 2762
rect 5017 2691 5070 2728
rect 5124 2754 5177 2838
rect 5124 2720 5132 2754
rect 5166 2720 5177 2754
rect 4960 2660 4972 2691
rect 5124 2690 5177 2720
rect 5207 2826 5261 2838
rect 5207 2792 5218 2826
rect 5252 2792 5261 2826
rect 5207 2736 5261 2792
rect 5207 2702 5218 2736
rect 5252 2702 5261 2736
rect 5207 2690 5261 2702
rect 5661 2824 5718 2836
rect 5661 2790 5673 2824
rect 5707 2790 5718 2824
rect 5661 2734 5718 2790
rect 5661 2700 5673 2734
rect 5707 2700 5718 2734
rect 5661 2688 5718 2700
rect 5748 2817 5798 2836
rect 5748 2696 5841 2817
rect 5748 2688 5777 2696
rect 5763 2662 5777 2688
rect 5811 2689 5841 2696
rect 5871 2689 5919 2817
rect 5949 2689 5997 2817
rect 6027 2741 6105 2817
rect 6027 2707 6038 2741
rect 6072 2707 6105 2741
rect 6027 2689 6105 2707
rect 6135 2748 6207 2817
rect 6135 2714 6154 2748
rect 6188 2714 6207 2748
rect 6135 2689 6207 2714
rect 6237 2696 6325 2817
rect 6237 2689 6264 2696
rect 5811 2662 5826 2689
rect 4914 2652 4972 2660
rect 5763 2650 5826 2662
rect 6252 2662 6264 2689
rect 6298 2689 6325 2696
rect 6355 2748 6411 2817
rect 6355 2714 6366 2748
rect 6400 2714 6411 2748
rect 6355 2689 6411 2714
rect 6441 2740 6540 2817
rect 6441 2706 6480 2740
rect 6514 2706 6540 2740
rect 6441 2689 6540 2706
rect 6570 2689 6618 2817
rect 6648 2751 6704 2817
rect 6648 2717 6659 2751
rect 6693 2717 6704 2751
rect 6648 2689 6704 2717
rect 6734 2699 6916 2817
rect 6734 2689 6761 2699
rect 6298 2662 6310 2689
rect 6749 2665 6761 2689
rect 6795 2665 6855 2699
rect 6889 2689 6916 2699
rect 6946 2692 7061 2817
rect 6946 2689 7000 2692
rect 6889 2665 6901 2689
rect 6252 2650 6310 2662
rect 6749 2653 6901 2665
rect 6988 2658 7000 2689
rect 7034 2689 7061 2692
rect 7091 2760 7144 2817
rect 7091 2726 7102 2760
rect 7136 2726 7144 2760
rect 7091 2689 7144 2726
rect 7198 2752 7251 2836
rect 7198 2718 7206 2752
rect 7240 2718 7251 2752
rect 7034 2658 7046 2689
rect 7198 2688 7251 2718
rect 7281 2824 7335 2836
rect 7281 2790 7292 2824
rect 7326 2790 7335 2824
rect 7281 2734 7335 2790
rect 7281 2700 7292 2734
rect 7326 2700 7335 2734
rect 7281 2688 7335 2700
rect 7723 2820 7780 2832
rect 7723 2786 7735 2820
rect 7769 2786 7780 2820
rect 7723 2730 7780 2786
rect 7723 2696 7735 2730
rect 7769 2696 7780 2730
rect 7723 2684 7780 2696
rect 7810 2813 7860 2832
rect 7810 2692 7903 2813
rect 7810 2684 7839 2692
rect 7825 2658 7839 2684
rect 7873 2685 7903 2692
rect 7933 2685 7981 2813
rect 8011 2685 8059 2813
rect 8089 2737 8167 2813
rect 8089 2703 8100 2737
rect 8134 2703 8167 2737
rect 8089 2685 8167 2703
rect 8197 2744 8269 2813
rect 8197 2710 8216 2744
rect 8250 2710 8269 2744
rect 8197 2685 8269 2710
rect 8299 2692 8387 2813
rect 8299 2685 8326 2692
rect 7873 2658 7888 2685
rect 6988 2650 7046 2658
rect 7825 2646 7888 2658
rect 8314 2658 8326 2685
rect 8360 2685 8387 2692
rect 8417 2744 8473 2813
rect 8417 2710 8428 2744
rect 8462 2710 8473 2744
rect 8417 2685 8473 2710
rect 8503 2736 8602 2813
rect 8503 2702 8542 2736
rect 8576 2702 8602 2736
rect 8503 2685 8602 2702
rect 8632 2685 8680 2813
rect 8710 2747 8766 2813
rect 8710 2713 8721 2747
rect 8755 2713 8766 2747
rect 8710 2685 8766 2713
rect 8796 2695 8978 2813
rect 8796 2685 8823 2695
rect 8360 2658 8372 2685
rect 8811 2661 8823 2685
rect 8857 2661 8917 2695
rect 8951 2685 8978 2695
rect 9008 2688 9123 2813
rect 9008 2685 9062 2688
rect 8951 2661 8963 2685
rect 8314 2646 8372 2658
rect 8811 2649 8963 2661
rect 9050 2654 9062 2685
rect 9096 2685 9123 2688
rect 9153 2756 9206 2813
rect 9153 2722 9164 2756
rect 9198 2722 9206 2756
rect 9153 2685 9206 2722
rect 9260 2748 9313 2832
rect 9260 2714 9268 2748
rect 9302 2714 9313 2748
rect 9096 2654 9108 2685
rect 9260 2684 9313 2714
rect 9343 2820 9397 2832
rect 9343 2786 9354 2820
rect 9388 2786 9397 2820
rect 9343 2730 9397 2786
rect 9343 2696 9354 2730
rect 9388 2696 9397 2730
rect 9343 2684 9397 2696
rect 9783 2816 9840 2828
rect 9783 2782 9795 2816
rect 9829 2782 9840 2816
rect 9783 2726 9840 2782
rect 9783 2692 9795 2726
rect 9829 2692 9840 2726
rect 9783 2680 9840 2692
rect 9870 2809 9920 2828
rect 9870 2688 9963 2809
rect 9870 2680 9899 2688
rect 9885 2654 9899 2680
rect 9933 2681 9963 2688
rect 9993 2681 10041 2809
rect 10071 2681 10119 2809
rect 10149 2733 10227 2809
rect 10149 2699 10160 2733
rect 10194 2699 10227 2733
rect 10149 2681 10227 2699
rect 10257 2740 10329 2809
rect 10257 2706 10276 2740
rect 10310 2706 10329 2740
rect 10257 2681 10329 2706
rect 10359 2688 10447 2809
rect 10359 2681 10386 2688
rect 9933 2654 9948 2681
rect 9050 2646 9108 2654
rect 9885 2642 9948 2654
rect 10374 2654 10386 2681
rect 10420 2681 10447 2688
rect 10477 2740 10533 2809
rect 10477 2706 10488 2740
rect 10522 2706 10533 2740
rect 10477 2681 10533 2706
rect 10563 2732 10662 2809
rect 10563 2698 10602 2732
rect 10636 2698 10662 2732
rect 10563 2681 10662 2698
rect 10692 2681 10740 2809
rect 10770 2743 10826 2809
rect 10770 2709 10781 2743
rect 10815 2709 10826 2743
rect 10770 2681 10826 2709
rect 10856 2691 11038 2809
rect 10856 2681 10883 2691
rect 10420 2654 10432 2681
rect 10871 2657 10883 2681
rect 10917 2657 10977 2691
rect 11011 2681 11038 2691
rect 11068 2684 11183 2809
rect 11068 2681 11122 2684
rect 11011 2657 11023 2681
rect 10374 2642 10432 2654
rect 10871 2645 11023 2657
rect 11110 2650 11122 2681
rect 11156 2681 11183 2684
rect 11213 2752 11266 2809
rect 11213 2718 11224 2752
rect 11258 2718 11266 2752
rect 11213 2681 11266 2718
rect 11320 2744 11373 2828
rect 11320 2710 11328 2744
rect 11362 2710 11373 2744
rect 11156 2650 11168 2681
rect 11320 2680 11373 2710
rect 11403 2816 11457 2828
rect 11403 2782 11414 2816
rect 11448 2782 11457 2816
rect 11403 2726 11457 2782
rect 11403 2692 11414 2726
rect 11448 2692 11457 2726
rect 11403 2680 11457 2692
rect 11845 2812 11902 2824
rect 11845 2778 11857 2812
rect 11891 2778 11902 2812
rect 11845 2722 11902 2778
rect 11845 2688 11857 2722
rect 11891 2688 11902 2722
rect 11845 2676 11902 2688
rect 11932 2805 11982 2824
rect 11932 2684 12025 2805
rect 11932 2676 11961 2684
rect 11947 2650 11961 2676
rect 11995 2677 12025 2684
rect 12055 2677 12103 2805
rect 12133 2677 12181 2805
rect 12211 2729 12289 2805
rect 12211 2695 12222 2729
rect 12256 2695 12289 2729
rect 12211 2677 12289 2695
rect 12319 2736 12391 2805
rect 12319 2702 12338 2736
rect 12372 2702 12391 2736
rect 12319 2677 12391 2702
rect 12421 2684 12509 2805
rect 12421 2677 12448 2684
rect 11995 2650 12010 2677
rect 11110 2642 11168 2650
rect 11947 2638 12010 2650
rect 12436 2650 12448 2677
rect 12482 2677 12509 2684
rect 12539 2736 12595 2805
rect 12539 2702 12550 2736
rect 12584 2702 12595 2736
rect 12539 2677 12595 2702
rect 12625 2728 12724 2805
rect 12625 2694 12664 2728
rect 12698 2694 12724 2728
rect 12625 2677 12724 2694
rect 12754 2677 12802 2805
rect 12832 2739 12888 2805
rect 12832 2705 12843 2739
rect 12877 2705 12888 2739
rect 12832 2677 12888 2705
rect 12918 2687 13100 2805
rect 12918 2677 12945 2687
rect 12482 2650 12494 2677
rect 12933 2653 12945 2677
rect 12979 2653 13039 2687
rect 13073 2677 13100 2687
rect 13130 2680 13245 2805
rect 13130 2677 13184 2680
rect 13073 2653 13085 2677
rect 12436 2638 12494 2650
rect 12933 2641 13085 2653
rect 13172 2646 13184 2677
rect 13218 2677 13245 2680
rect 13275 2748 13328 2805
rect 13275 2714 13286 2748
rect 13320 2714 13328 2748
rect 13275 2677 13328 2714
rect 13382 2740 13435 2824
rect 13382 2706 13390 2740
rect 13424 2706 13435 2740
rect 13218 2646 13230 2677
rect 13382 2676 13435 2706
rect 13465 2812 13519 2824
rect 13465 2778 13476 2812
rect 13510 2778 13519 2812
rect 13465 2722 13519 2778
rect 13465 2688 13476 2722
rect 13510 2688 13519 2722
rect 13465 2676 13519 2688
rect 13919 2810 13976 2822
rect 13919 2776 13931 2810
rect 13965 2776 13976 2810
rect 13919 2720 13976 2776
rect 13919 2686 13931 2720
rect 13965 2686 13976 2720
rect 13919 2674 13976 2686
rect 14006 2803 14056 2822
rect 14006 2682 14099 2803
rect 14006 2674 14035 2682
rect 14021 2648 14035 2674
rect 14069 2675 14099 2682
rect 14129 2675 14177 2803
rect 14207 2675 14255 2803
rect 14285 2727 14363 2803
rect 14285 2693 14296 2727
rect 14330 2693 14363 2727
rect 14285 2675 14363 2693
rect 14393 2734 14465 2803
rect 14393 2700 14412 2734
rect 14446 2700 14465 2734
rect 14393 2675 14465 2700
rect 14495 2682 14583 2803
rect 14495 2675 14522 2682
rect 14069 2648 14084 2675
rect 13172 2638 13230 2646
rect 14021 2636 14084 2648
rect 14510 2648 14522 2675
rect 14556 2675 14583 2682
rect 14613 2734 14669 2803
rect 14613 2700 14624 2734
rect 14658 2700 14669 2734
rect 14613 2675 14669 2700
rect 14699 2726 14798 2803
rect 14699 2692 14738 2726
rect 14772 2692 14798 2726
rect 14699 2675 14798 2692
rect 14828 2675 14876 2803
rect 14906 2737 14962 2803
rect 14906 2703 14917 2737
rect 14951 2703 14962 2737
rect 14906 2675 14962 2703
rect 14992 2685 15174 2803
rect 14992 2675 15019 2685
rect 14556 2648 14568 2675
rect 15007 2651 15019 2675
rect 15053 2651 15113 2685
rect 15147 2675 15174 2685
rect 15204 2678 15319 2803
rect 15204 2675 15258 2678
rect 15147 2651 15159 2675
rect 14510 2636 14568 2648
rect 15007 2639 15159 2651
rect 15246 2644 15258 2675
rect 15292 2675 15319 2678
rect 15349 2746 15402 2803
rect 15349 2712 15360 2746
rect 15394 2712 15402 2746
rect 15349 2675 15402 2712
rect 15456 2738 15509 2822
rect 15456 2704 15464 2738
rect 15498 2704 15509 2738
rect 15292 2644 15304 2675
rect 15456 2674 15509 2704
rect 15539 2810 15593 2822
rect 15539 2776 15550 2810
rect 15584 2776 15593 2810
rect 15539 2720 15593 2776
rect 15539 2686 15550 2720
rect 15584 2686 15593 2720
rect 15539 2674 15593 2686
rect 15981 2806 16038 2818
rect 15981 2772 15993 2806
rect 16027 2772 16038 2806
rect 15981 2716 16038 2772
rect 15981 2682 15993 2716
rect 16027 2682 16038 2716
rect 15981 2670 16038 2682
rect 16068 2799 16118 2818
rect 16068 2678 16161 2799
rect 16068 2670 16097 2678
rect 16083 2644 16097 2670
rect 16131 2671 16161 2678
rect 16191 2671 16239 2799
rect 16269 2671 16317 2799
rect 16347 2723 16425 2799
rect 16347 2689 16358 2723
rect 16392 2689 16425 2723
rect 16347 2671 16425 2689
rect 16455 2730 16527 2799
rect 16455 2696 16474 2730
rect 16508 2696 16527 2730
rect 16455 2671 16527 2696
rect 16557 2678 16645 2799
rect 16557 2671 16584 2678
rect 16131 2644 16146 2671
rect 15246 2636 15304 2644
rect 16083 2632 16146 2644
rect 16572 2644 16584 2671
rect 16618 2671 16645 2678
rect 16675 2730 16731 2799
rect 16675 2696 16686 2730
rect 16720 2696 16731 2730
rect 16675 2671 16731 2696
rect 16761 2722 16860 2799
rect 16761 2688 16800 2722
rect 16834 2688 16860 2722
rect 16761 2671 16860 2688
rect 16890 2671 16938 2799
rect 16968 2733 17024 2799
rect 16968 2699 16979 2733
rect 17013 2699 17024 2733
rect 16968 2671 17024 2699
rect 17054 2681 17236 2799
rect 17054 2671 17081 2681
rect 16618 2644 16630 2671
rect 17069 2647 17081 2671
rect 17115 2647 17175 2681
rect 17209 2671 17236 2681
rect 17266 2674 17381 2799
rect 17266 2671 17320 2674
rect 17209 2647 17221 2671
rect 16572 2632 16630 2644
rect 17069 2635 17221 2647
rect 17308 2640 17320 2671
rect 17354 2671 17381 2674
rect 17411 2742 17464 2799
rect 17411 2708 17422 2742
rect 17456 2708 17464 2742
rect 17411 2671 17464 2708
rect 17518 2734 17571 2818
rect 17518 2700 17526 2734
rect 17560 2700 17571 2734
rect 17354 2640 17366 2671
rect 17518 2670 17571 2700
rect 17601 2806 17655 2818
rect 17601 2772 17612 2806
rect 17646 2772 17655 2806
rect 17601 2716 17655 2772
rect 17601 2682 17612 2716
rect 17646 2682 17655 2716
rect 17601 2670 17655 2682
rect 17308 2632 17366 2640
<< pdiff >>
rect 18190 6085 18242 6097
rect 18190 6051 18198 6085
rect 18232 6051 18242 6085
rect 18190 6017 18242 6051
rect 18190 5983 18198 6017
rect 18232 5983 18242 6017
rect 18190 5949 18242 5983
rect 18190 5915 18198 5949
rect 18232 5915 18242 5949
rect 18190 5897 18242 5915
rect 18272 6085 18324 6097
rect 18272 6051 18282 6085
rect 18316 6051 18324 6085
rect 18272 6017 18324 6051
rect 18272 5983 18282 6017
rect 18316 5983 18324 6017
rect 18272 5949 18324 5983
rect 18272 5915 18282 5949
rect 18316 5915 18324 5949
rect 18272 5897 18324 5915
rect 26332 6037 26384 6049
rect 26332 6003 26340 6037
rect 26374 6003 26384 6037
rect 26332 5969 26384 6003
rect 26332 5935 26340 5969
rect 26374 5935 26384 5969
rect 26332 5899 26384 5935
rect 26332 5865 26340 5899
rect 26374 5865 26384 5899
rect 26332 5849 26384 5865
rect 26414 6037 26468 6049
rect 26414 6003 26424 6037
rect 26458 6003 26468 6037
rect 26414 5969 26468 6003
rect 26414 5935 26424 5969
rect 26458 5935 26468 5969
rect 26414 5899 26468 5935
rect 26414 5865 26424 5899
rect 26458 5865 26468 5899
rect 26414 5849 26468 5865
rect 26498 6037 26552 6049
rect 26498 6003 26508 6037
rect 26542 6003 26552 6037
rect 26498 5969 26552 6003
rect 26498 5935 26508 5969
rect 26542 5935 26552 5969
rect 26498 5849 26552 5935
rect 26582 6037 26636 6049
rect 26582 6003 26592 6037
rect 26626 6003 26636 6037
rect 26582 5969 26636 6003
rect 26582 5935 26592 5969
rect 26626 5935 26636 5969
rect 26582 5899 26636 5935
rect 26582 5865 26592 5899
rect 26626 5865 26636 5899
rect 26582 5849 26636 5865
rect 26666 6037 26720 6049
rect 26666 6003 26676 6037
rect 26710 6003 26720 6037
rect 26666 5969 26720 6003
rect 26666 5935 26676 5969
rect 26710 5935 26720 5969
rect 26666 5849 26720 5935
rect 26750 6037 26804 6049
rect 26750 6003 26760 6037
rect 26794 6003 26804 6037
rect 26750 5969 26804 6003
rect 26750 5935 26760 5969
rect 26794 5935 26804 5969
rect 26750 5899 26804 5935
rect 26750 5865 26760 5899
rect 26794 5865 26804 5899
rect 26750 5849 26804 5865
rect 26834 6037 26888 6049
rect 26834 6003 26844 6037
rect 26878 6003 26888 6037
rect 26834 5969 26888 6003
rect 26834 5935 26844 5969
rect 26878 5935 26888 5969
rect 26834 5849 26888 5935
rect 26918 6037 26972 6049
rect 26918 6003 26928 6037
rect 26962 6003 26972 6037
rect 26918 5969 26972 6003
rect 26918 5935 26928 5969
rect 26962 5935 26972 5969
rect 26918 5899 26972 5935
rect 26918 5865 26928 5899
rect 26962 5865 26972 5899
rect 26918 5849 26972 5865
rect 27002 6037 27056 6049
rect 27002 6003 27012 6037
rect 27046 6003 27056 6037
rect 27002 5969 27056 6003
rect 27002 5935 27012 5969
rect 27046 5935 27056 5969
rect 27002 5849 27056 5935
rect 27086 6037 27140 6049
rect 27086 6003 27096 6037
rect 27130 6003 27140 6037
rect 27086 5969 27140 6003
rect 27086 5935 27096 5969
rect 27130 5935 27140 5969
rect 27086 5899 27140 5935
rect 27086 5865 27096 5899
rect 27130 5865 27140 5899
rect 27086 5849 27140 5865
rect 27170 6037 27224 6049
rect 27170 6003 27180 6037
rect 27214 6003 27224 6037
rect 27170 5969 27224 6003
rect 27170 5935 27180 5969
rect 27214 5935 27224 5969
rect 27170 5849 27224 5935
rect 27254 6037 27308 6049
rect 27254 6003 27264 6037
rect 27298 6003 27308 6037
rect 27254 5969 27308 6003
rect 27254 5935 27264 5969
rect 27298 5935 27308 5969
rect 27254 5899 27308 5935
rect 27254 5865 27264 5899
rect 27298 5865 27308 5899
rect 27254 5849 27308 5865
rect 27338 6037 27392 6049
rect 27338 6003 27348 6037
rect 27382 6003 27392 6037
rect 27338 5969 27392 6003
rect 27338 5935 27348 5969
rect 27382 5935 27392 5969
rect 27338 5849 27392 5935
rect 27422 6037 27476 6049
rect 27422 6003 27432 6037
rect 27466 6003 27476 6037
rect 27422 5969 27476 6003
rect 27422 5935 27432 5969
rect 27466 5935 27476 5969
rect 27422 5899 27476 5935
rect 27422 5865 27432 5899
rect 27466 5865 27476 5899
rect 27422 5849 27476 5865
rect 27506 6037 27560 6049
rect 27506 6003 27516 6037
rect 27550 6003 27560 6037
rect 27506 5969 27560 6003
rect 27506 5935 27516 5969
rect 27550 5935 27560 5969
rect 27506 5849 27560 5935
rect 27590 6037 27644 6049
rect 27590 6003 27600 6037
rect 27634 6003 27644 6037
rect 27590 5969 27644 6003
rect 27590 5935 27600 5969
rect 27634 5935 27644 5969
rect 27590 5899 27644 5935
rect 27590 5865 27600 5899
rect 27634 5865 27644 5899
rect 27590 5849 27644 5865
rect 27674 6037 27726 6049
rect 27674 6003 27684 6037
rect 27718 6003 27726 6037
rect 27674 5969 27726 6003
rect 27674 5935 27684 5969
rect 27718 5935 27726 5969
rect 27674 5849 27726 5935
rect 28138 6019 28190 6031
rect 28138 5985 28146 6019
rect 28180 5985 28190 6019
rect 28138 5951 28190 5985
rect 28138 5917 28146 5951
rect 28180 5917 28190 5951
rect 28138 5881 28190 5917
rect 28138 5847 28146 5881
rect 28180 5847 28190 5881
rect 28138 5831 28190 5847
rect 28220 6019 28274 6031
rect 28220 5985 28230 6019
rect 28264 5985 28274 6019
rect 28220 5951 28274 5985
rect 28220 5917 28230 5951
rect 28264 5917 28274 5951
rect 28220 5881 28274 5917
rect 28220 5847 28230 5881
rect 28264 5847 28274 5881
rect 28220 5831 28274 5847
rect 28304 6019 28358 6031
rect 28304 5985 28314 6019
rect 28348 5985 28358 6019
rect 28304 5951 28358 5985
rect 28304 5917 28314 5951
rect 28348 5917 28358 5951
rect 28304 5831 28358 5917
rect 28388 6019 28442 6031
rect 28388 5985 28398 6019
rect 28432 5985 28442 6019
rect 28388 5951 28442 5985
rect 28388 5917 28398 5951
rect 28432 5917 28442 5951
rect 28388 5881 28442 5917
rect 28388 5847 28398 5881
rect 28432 5847 28442 5881
rect 28388 5831 28442 5847
rect 28472 6019 28526 6031
rect 28472 5985 28482 6019
rect 28516 5985 28526 6019
rect 28472 5951 28526 5985
rect 28472 5917 28482 5951
rect 28516 5917 28526 5951
rect 28472 5831 28526 5917
rect 28556 6019 28610 6031
rect 28556 5985 28566 6019
rect 28600 5985 28610 6019
rect 28556 5951 28610 5985
rect 28556 5917 28566 5951
rect 28600 5917 28610 5951
rect 28556 5881 28610 5917
rect 28556 5847 28566 5881
rect 28600 5847 28610 5881
rect 28556 5831 28610 5847
rect 28640 6019 28694 6031
rect 28640 5985 28650 6019
rect 28684 5985 28694 6019
rect 28640 5951 28694 5985
rect 28640 5917 28650 5951
rect 28684 5917 28694 5951
rect 28640 5831 28694 5917
rect 28724 6019 28778 6031
rect 28724 5985 28734 6019
rect 28768 5985 28778 6019
rect 28724 5951 28778 5985
rect 28724 5917 28734 5951
rect 28768 5917 28778 5951
rect 28724 5881 28778 5917
rect 28724 5847 28734 5881
rect 28768 5847 28778 5881
rect 28724 5831 28778 5847
rect 28808 6019 28862 6031
rect 28808 5985 28818 6019
rect 28852 5985 28862 6019
rect 28808 5951 28862 5985
rect 28808 5917 28818 5951
rect 28852 5917 28862 5951
rect 28808 5831 28862 5917
rect 28892 6019 28946 6031
rect 28892 5985 28902 6019
rect 28936 5985 28946 6019
rect 28892 5951 28946 5985
rect 28892 5917 28902 5951
rect 28936 5917 28946 5951
rect 28892 5881 28946 5917
rect 28892 5847 28902 5881
rect 28936 5847 28946 5881
rect 28892 5831 28946 5847
rect 28976 6019 29030 6031
rect 28976 5985 28986 6019
rect 29020 5985 29030 6019
rect 28976 5951 29030 5985
rect 28976 5917 28986 5951
rect 29020 5917 29030 5951
rect 28976 5831 29030 5917
rect 29060 6019 29114 6031
rect 29060 5985 29070 6019
rect 29104 5985 29114 6019
rect 29060 5951 29114 5985
rect 29060 5917 29070 5951
rect 29104 5917 29114 5951
rect 29060 5881 29114 5917
rect 29060 5847 29070 5881
rect 29104 5847 29114 5881
rect 29060 5831 29114 5847
rect 29144 6019 29198 6031
rect 29144 5985 29154 6019
rect 29188 5985 29198 6019
rect 29144 5951 29198 5985
rect 29144 5917 29154 5951
rect 29188 5917 29198 5951
rect 29144 5831 29198 5917
rect 29228 6019 29282 6031
rect 29228 5985 29238 6019
rect 29272 5985 29282 6019
rect 29228 5951 29282 5985
rect 29228 5917 29238 5951
rect 29272 5917 29282 5951
rect 29228 5881 29282 5917
rect 29228 5847 29238 5881
rect 29272 5847 29282 5881
rect 29228 5831 29282 5847
rect 29312 6019 29366 6031
rect 29312 5985 29322 6019
rect 29356 5985 29366 6019
rect 29312 5951 29366 5985
rect 29312 5917 29322 5951
rect 29356 5917 29366 5951
rect 29312 5831 29366 5917
rect 29396 6019 29450 6031
rect 29396 5985 29406 6019
rect 29440 5985 29450 6019
rect 29396 5951 29450 5985
rect 29396 5917 29406 5951
rect 29440 5917 29450 5951
rect 29396 5881 29450 5917
rect 29396 5847 29406 5881
rect 29440 5847 29450 5881
rect 29396 5831 29450 5847
rect 29480 6019 29532 6031
rect 29480 5985 29490 6019
rect 29524 5985 29532 6019
rect 29480 5951 29532 5985
rect 29480 5917 29490 5951
rect 29524 5917 29532 5951
rect 29480 5831 29532 5917
rect 1525 3200 1582 3212
rect 1525 3166 1535 3200
rect 1569 3166 1582 3200
rect 1525 3117 1582 3166
rect 1525 3083 1535 3117
rect 1569 3083 1582 3117
rect 1525 3034 1582 3083
rect 1525 3000 1535 3034
rect 1569 3000 1582 3034
rect 1525 2988 1582 3000
rect 1612 3200 1667 3212
rect 1612 3166 1625 3200
rect 1659 3188 1667 3200
rect 1733 3188 1786 3209
rect 1659 3166 1685 3188
rect 1612 3132 1685 3166
rect 1612 3098 1625 3132
rect 1659 3098 1685 3132
rect 1612 3064 1685 3098
rect 1612 3030 1625 3064
rect 1659 3030 1685 3064
rect 1612 2988 1685 3030
rect 1715 3009 1786 3188
rect 1816 3167 1869 3209
rect 2122 3196 2173 3208
rect 2122 3167 2130 3196
rect 1816 3009 1887 3167
rect 1715 2988 1768 3009
rect 1834 2967 1887 3009
rect 1917 3155 1977 3167
rect 1917 3121 1930 3155
rect 1964 3121 1977 3155
rect 1917 3087 1977 3121
rect 1917 3053 1930 3087
rect 1964 3053 1977 3087
rect 1917 3019 1977 3053
rect 1917 2985 1930 3019
rect 1964 2985 1977 3019
rect 1917 2967 1977 2985
rect 2007 3155 2074 3167
rect 2007 3121 2020 3155
rect 2054 3121 2074 3155
rect 2007 3063 2074 3121
rect 2007 3029 2020 3063
rect 2054 3029 2074 3063
rect 2007 2967 2074 3029
rect 2104 3162 2130 3167
rect 2164 3167 2173 3196
rect 3053 3200 3112 3212
rect 2742 3167 2861 3182
rect 2164 3162 2191 3167
rect 2104 2967 2191 3162
rect 2221 3128 2292 3167
rect 2221 3094 2234 3128
rect 2268 3094 2292 3128
rect 2221 2967 2292 3094
rect 2322 3131 2384 3167
rect 2322 3097 2335 3131
rect 2369 3097 2384 3131
rect 2322 2967 2384 3097
rect 2414 2967 2485 3167
rect 2515 3155 2575 3167
rect 2515 3121 2528 3155
rect 2562 3121 2575 3155
rect 2515 3044 2575 3121
rect 2515 3010 2528 3044
rect 2562 3010 2575 3044
rect 2515 2967 2575 3010
rect 2605 3155 2694 3167
rect 2605 3121 2647 3155
rect 2681 3121 2694 3155
rect 2605 3071 2694 3121
rect 2605 3037 2647 3071
rect 2681 3037 2694 3071
rect 2605 2967 2694 3037
rect 2724 3157 2861 3167
rect 2724 3123 2738 3157
rect 2772 3123 2813 3157
rect 2847 3123 2861 3157
rect 2724 2982 2861 3123
rect 2891 3170 2958 3182
rect 2891 3136 2912 3170
rect 2946 3136 2958 3170
rect 2891 3060 2958 3136
rect 2891 3026 2912 3060
rect 2946 3026 2958 3060
rect 2891 2982 2958 3026
rect 3053 3166 3065 3200
rect 3099 3166 3112 3200
rect 3053 3117 3112 3166
rect 3053 3083 3065 3117
rect 3099 3083 3112 3117
rect 3053 3034 3112 3083
rect 3053 3000 3065 3034
rect 3099 3000 3112 3034
rect 3053 2988 3112 3000
rect 3142 3200 3199 3212
rect 3142 3166 3155 3200
rect 3189 3166 3199 3200
rect 3142 3117 3199 3166
rect 3142 3083 3155 3117
rect 3189 3083 3199 3117
rect 3142 3034 3199 3083
rect 3142 3000 3155 3034
rect 3189 3000 3199 3034
rect 3142 2988 3199 3000
rect 3587 3196 3644 3208
rect 3587 3162 3597 3196
rect 3631 3162 3644 3196
rect 3587 3113 3644 3162
rect 3587 3079 3597 3113
rect 3631 3079 3644 3113
rect 3587 3030 3644 3079
rect 3587 2996 3597 3030
rect 3631 2996 3644 3030
rect 2724 2967 2777 2982
rect 3587 2984 3644 2996
rect 3674 3196 3729 3208
rect 3674 3162 3687 3196
rect 3721 3184 3729 3196
rect 3795 3184 3848 3205
rect 3721 3162 3747 3184
rect 3674 3128 3747 3162
rect 3674 3094 3687 3128
rect 3721 3094 3747 3128
rect 3674 3060 3747 3094
rect 3674 3026 3687 3060
rect 3721 3026 3747 3060
rect 3674 2984 3747 3026
rect 3777 3005 3848 3184
rect 3878 3163 3931 3205
rect 4184 3192 4235 3204
rect 4184 3163 4192 3192
rect 3878 3005 3949 3163
rect 3777 2984 3830 3005
rect 3896 2963 3949 3005
rect 3979 3151 4039 3163
rect 3979 3117 3992 3151
rect 4026 3117 4039 3151
rect 3979 3083 4039 3117
rect 3979 3049 3992 3083
rect 4026 3049 4039 3083
rect 3979 3015 4039 3049
rect 3979 2981 3992 3015
rect 4026 2981 4039 3015
rect 3979 2963 4039 2981
rect 4069 3151 4136 3163
rect 4069 3117 4082 3151
rect 4116 3117 4136 3151
rect 4069 3059 4136 3117
rect 4069 3025 4082 3059
rect 4116 3025 4136 3059
rect 4069 2963 4136 3025
rect 4166 3158 4192 3163
rect 4226 3163 4235 3192
rect 5115 3196 5174 3208
rect 4804 3163 4923 3178
rect 4226 3158 4253 3163
rect 4166 2963 4253 3158
rect 4283 3124 4354 3163
rect 4283 3090 4296 3124
rect 4330 3090 4354 3124
rect 4283 2963 4354 3090
rect 4384 3127 4446 3163
rect 4384 3093 4397 3127
rect 4431 3093 4446 3127
rect 4384 2963 4446 3093
rect 4476 2963 4547 3163
rect 4577 3151 4637 3163
rect 4577 3117 4590 3151
rect 4624 3117 4637 3151
rect 4577 3040 4637 3117
rect 4577 3006 4590 3040
rect 4624 3006 4637 3040
rect 4577 2963 4637 3006
rect 4667 3151 4756 3163
rect 4667 3117 4709 3151
rect 4743 3117 4756 3151
rect 4667 3067 4756 3117
rect 4667 3033 4709 3067
rect 4743 3033 4756 3067
rect 4667 2963 4756 3033
rect 4786 3153 4923 3163
rect 4786 3119 4800 3153
rect 4834 3119 4875 3153
rect 4909 3119 4923 3153
rect 4786 2978 4923 3119
rect 4953 3166 5020 3178
rect 4953 3132 4974 3166
rect 5008 3132 5020 3166
rect 4953 3056 5020 3132
rect 4953 3022 4974 3056
rect 5008 3022 5020 3056
rect 4953 2978 5020 3022
rect 5115 3162 5127 3196
rect 5161 3162 5174 3196
rect 5115 3113 5174 3162
rect 5115 3079 5127 3113
rect 5161 3079 5174 3113
rect 5115 3030 5174 3079
rect 5115 2996 5127 3030
rect 5161 2996 5174 3030
rect 5115 2984 5174 2996
rect 5204 3196 5261 3208
rect 5204 3162 5217 3196
rect 5251 3162 5261 3196
rect 5204 3113 5261 3162
rect 5204 3079 5217 3113
rect 5251 3079 5261 3113
rect 5204 3030 5261 3079
rect 5204 2996 5217 3030
rect 5251 2996 5261 3030
rect 5204 2984 5261 2996
rect 5661 3194 5718 3206
rect 5661 3160 5671 3194
rect 5705 3160 5718 3194
rect 5661 3111 5718 3160
rect 5661 3077 5671 3111
rect 5705 3077 5718 3111
rect 5661 3028 5718 3077
rect 5661 2994 5671 3028
rect 5705 2994 5718 3028
rect 4786 2963 4839 2978
rect 5661 2982 5718 2994
rect 5748 3194 5803 3206
rect 5748 3160 5761 3194
rect 5795 3182 5803 3194
rect 5869 3182 5922 3203
rect 5795 3160 5821 3182
rect 5748 3126 5821 3160
rect 5748 3092 5761 3126
rect 5795 3092 5821 3126
rect 5748 3058 5821 3092
rect 5748 3024 5761 3058
rect 5795 3024 5821 3058
rect 5748 2982 5821 3024
rect 5851 3003 5922 3182
rect 5952 3161 6005 3203
rect 6258 3190 6309 3202
rect 6258 3161 6266 3190
rect 5952 3003 6023 3161
rect 5851 2982 5904 3003
rect 5970 2961 6023 3003
rect 6053 3149 6113 3161
rect 6053 3115 6066 3149
rect 6100 3115 6113 3149
rect 6053 3081 6113 3115
rect 6053 3047 6066 3081
rect 6100 3047 6113 3081
rect 6053 3013 6113 3047
rect 6053 2979 6066 3013
rect 6100 2979 6113 3013
rect 6053 2961 6113 2979
rect 6143 3149 6210 3161
rect 6143 3115 6156 3149
rect 6190 3115 6210 3149
rect 6143 3057 6210 3115
rect 6143 3023 6156 3057
rect 6190 3023 6210 3057
rect 6143 2961 6210 3023
rect 6240 3156 6266 3161
rect 6300 3161 6309 3190
rect 7189 3194 7248 3206
rect 6878 3161 6997 3176
rect 6300 3156 6327 3161
rect 6240 2961 6327 3156
rect 6357 3122 6428 3161
rect 6357 3088 6370 3122
rect 6404 3088 6428 3122
rect 6357 2961 6428 3088
rect 6458 3125 6520 3161
rect 6458 3091 6471 3125
rect 6505 3091 6520 3125
rect 6458 2961 6520 3091
rect 6550 2961 6621 3161
rect 6651 3149 6711 3161
rect 6651 3115 6664 3149
rect 6698 3115 6711 3149
rect 6651 3038 6711 3115
rect 6651 3004 6664 3038
rect 6698 3004 6711 3038
rect 6651 2961 6711 3004
rect 6741 3149 6830 3161
rect 6741 3115 6783 3149
rect 6817 3115 6830 3149
rect 6741 3065 6830 3115
rect 6741 3031 6783 3065
rect 6817 3031 6830 3065
rect 6741 2961 6830 3031
rect 6860 3151 6997 3161
rect 6860 3117 6874 3151
rect 6908 3117 6949 3151
rect 6983 3117 6997 3151
rect 6860 2976 6997 3117
rect 7027 3164 7094 3176
rect 7027 3130 7048 3164
rect 7082 3130 7094 3164
rect 7027 3054 7094 3130
rect 7027 3020 7048 3054
rect 7082 3020 7094 3054
rect 7027 2976 7094 3020
rect 7189 3160 7201 3194
rect 7235 3160 7248 3194
rect 7189 3111 7248 3160
rect 7189 3077 7201 3111
rect 7235 3077 7248 3111
rect 7189 3028 7248 3077
rect 7189 2994 7201 3028
rect 7235 2994 7248 3028
rect 7189 2982 7248 2994
rect 7278 3194 7335 3206
rect 7278 3160 7291 3194
rect 7325 3160 7335 3194
rect 7278 3111 7335 3160
rect 7278 3077 7291 3111
rect 7325 3077 7335 3111
rect 7278 3028 7335 3077
rect 7278 2994 7291 3028
rect 7325 2994 7335 3028
rect 7278 2982 7335 2994
rect 7723 3190 7780 3202
rect 7723 3156 7733 3190
rect 7767 3156 7780 3190
rect 7723 3107 7780 3156
rect 7723 3073 7733 3107
rect 7767 3073 7780 3107
rect 7723 3024 7780 3073
rect 7723 2990 7733 3024
rect 7767 2990 7780 3024
rect 6860 2961 6913 2976
rect 7723 2978 7780 2990
rect 7810 3190 7865 3202
rect 7810 3156 7823 3190
rect 7857 3178 7865 3190
rect 7931 3178 7984 3199
rect 7857 3156 7883 3178
rect 7810 3122 7883 3156
rect 7810 3088 7823 3122
rect 7857 3088 7883 3122
rect 7810 3054 7883 3088
rect 7810 3020 7823 3054
rect 7857 3020 7883 3054
rect 7810 2978 7883 3020
rect 7913 2999 7984 3178
rect 8014 3157 8067 3199
rect 8320 3186 8371 3198
rect 8320 3157 8328 3186
rect 8014 2999 8085 3157
rect 7913 2978 7966 2999
rect 8032 2957 8085 2999
rect 8115 3145 8175 3157
rect 8115 3111 8128 3145
rect 8162 3111 8175 3145
rect 8115 3077 8175 3111
rect 8115 3043 8128 3077
rect 8162 3043 8175 3077
rect 8115 3009 8175 3043
rect 8115 2975 8128 3009
rect 8162 2975 8175 3009
rect 8115 2957 8175 2975
rect 8205 3145 8272 3157
rect 8205 3111 8218 3145
rect 8252 3111 8272 3145
rect 8205 3053 8272 3111
rect 8205 3019 8218 3053
rect 8252 3019 8272 3053
rect 8205 2957 8272 3019
rect 8302 3152 8328 3157
rect 8362 3157 8371 3186
rect 9251 3190 9310 3202
rect 8940 3157 9059 3172
rect 8362 3152 8389 3157
rect 8302 2957 8389 3152
rect 8419 3118 8490 3157
rect 8419 3084 8432 3118
rect 8466 3084 8490 3118
rect 8419 2957 8490 3084
rect 8520 3121 8582 3157
rect 8520 3087 8533 3121
rect 8567 3087 8582 3121
rect 8520 2957 8582 3087
rect 8612 2957 8683 3157
rect 8713 3145 8773 3157
rect 8713 3111 8726 3145
rect 8760 3111 8773 3145
rect 8713 3034 8773 3111
rect 8713 3000 8726 3034
rect 8760 3000 8773 3034
rect 8713 2957 8773 3000
rect 8803 3145 8892 3157
rect 8803 3111 8845 3145
rect 8879 3111 8892 3145
rect 8803 3061 8892 3111
rect 8803 3027 8845 3061
rect 8879 3027 8892 3061
rect 8803 2957 8892 3027
rect 8922 3147 9059 3157
rect 8922 3113 8936 3147
rect 8970 3113 9011 3147
rect 9045 3113 9059 3147
rect 8922 2972 9059 3113
rect 9089 3160 9156 3172
rect 9089 3126 9110 3160
rect 9144 3126 9156 3160
rect 9089 3050 9156 3126
rect 9089 3016 9110 3050
rect 9144 3016 9156 3050
rect 9089 2972 9156 3016
rect 9251 3156 9263 3190
rect 9297 3156 9310 3190
rect 9251 3107 9310 3156
rect 9251 3073 9263 3107
rect 9297 3073 9310 3107
rect 9251 3024 9310 3073
rect 9251 2990 9263 3024
rect 9297 2990 9310 3024
rect 9251 2978 9310 2990
rect 9340 3190 9397 3202
rect 9340 3156 9353 3190
rect 9387 3156 9397 3190
rect 9340 3107 9397 3156
rect 9340 3073 9353 3107
rect 9387 3073 9397 3107
rect 9340 3024 9397 3073
rect 9340 2990 9353 3024
rect 9387 2990 9397 3024
rect 9340 2978 9397 2990
rect 9783 3186 9840 3198
rect 9783 3152 9793 3186
rect 9827 3152 9840 3186
rect 9783 3103 9840 3152
rect 9783 3069 9793 3103
rect 9827 3069 9840 3103
rect 9783 3020 9840 3069
rect 9783 2986 9793 3020
rect 9827 2986 9840 3020
rect 8922 2957 8975 2972
rect 9783 2974 9840 2986
rect 9870 3186 9925 3198
rect 9870 3152 9883 3186
rect 9917 3174 9925 3186
rect 9991 3174 10044 3195
rect 9917 3152 9943 3174
rect 9870 3118 9943 3152
rect 9870 3084 9883 3118
rect 9917 3084 9943 3118
rect 9870 3050 9943 3084
rect 9870 3016 9883 3050
rect 9917 3016 9943 3050
rect 9870 2974 9943 3016
rect 9973 2995 10044 3174
rect 10074 3153 10127 3195
rect 10380 3182 10431 3194
rect 10380 3153 10388 3182
rect 10074 2995 10145 3153
rect 9973 2974 10026 2995
rect 10092 2953 10145 2995
rect 10175 3141 10235 3153
rect 10175 3107 10188 3141
rect 10222 3107 10235 3141
rect 10175 3073 10235 3107
rect 10175 3039 10188 3073
rect 10222 3039 10235 3073
rect 10175 3005 10235 3039
rect 10175 2971 10188 3005
rect 10222 2971 10235 3005
rect 10175 2953 10235 2971
rect 10265 3141 10332 3153
rect 10265 3107 10278 3141
rect 10312 3107 10332 3141
rect 10265 3049 10332 3107
rect 10265 3015 10278 3049
rect 10312 3015 10332 3049
rect 10265 2953 10332 3015
rect 10362 3148 10388 3153
rect 10422 3153 10431 3182
rect 11311 3186 11370 3198
rect 11000 3153 11119 3168
rect 10422 3148 10449 3153
rect 10362 2953 10449 3148
rect 10479 3114 10550 3153
rect 10479 3080 10492 3114
rect 10526 3080 10550 3114
rect 10479 2953 10550 3080
rect 10580 3117 10642 3153
rect 10580 3083 10593 3117
rect 10627 3083 10642 3117
rect 10580 2953 10642 3083
rect 10672 2953 10743 3153
rect 10773 3141 10833 3153
rect 10773 3107 10786 3141
rect 10820 3107 10833 3141
rect 10773 3030 10833 3107
rect 10773 2996 10786 3030
rect 10820 2996 10833 3030
rect 10773 2953 10833 2996
rect 10863 3141 10952 3153
rect 10863 3107 10905 3141
rect 10939 3107 10952 3141
rect 10863 3057 10952 3107
rect 10863 3023 10905 3057
rect 10939 3023 10952 3057
rect 10863 2953 10952 3023
rect 10982 3143 11119 3153
rect 10982 3109 10996 3143
rect 11030 3109 11071 3143
rect 11105 3109 11119 3143
rect 10982 2968 11119 3109
rect 11149 3156 11216 3168
rect 11149 3122 11170 3156
rect 11204 3122 11216 3156
rect 11149 3046 11216 3122
rect 11149 3012 11170 3046
rect 11204 3012 11216 3046
rect 11149 2968 11216 3012
rect 11311 3152 11323 3186
rect 11357 3152 11370 3186
rect 11311 3103 11370 3152
rect 11311 3069 11323 3103
rect 11357 3069 11370 3103
rect 11311 3020 11370 3069
rect 11311 2986 11323 3020
rect 11357 2986 11370 3020
rect 11311 2974 11370 2986
rect 11400 3186 11457 3198
rect 11400 3152 11413 3186
rect 11447 3152 11457 3186
rect 11400 3103 11457 3152
rect 11400 3069 11413 3103
rect 11447 3069 11457 3103
rect 11400 3020 11457 3069
rect 11400 2986 11413 3020
rect 11447 2986 11457 3020
rect 11400 2974 11457 2986
rect 11845 3182 11902 3194
rect 11845 3148 11855 3182
rect 11889 3148 11902 3182
rect 11845 3099 11902 3148
rect 11845 3065 11855 3099
rect 11889 3065 11902 3099
rect 11845 3016 11902 3065
rect 11845 2982 11855 3016
rect 11889 2982 11902 3016
rect 10982 2953 11035 2968
rect 11845 2970 11902 2982
rect 11932 3182 11987 3194
rect 11932 3148 11945 3182
rect 11979 3170 11987 3182
rect 12053 3170 12106 3191
rect 11979 3148 12005 3170
rect 11932 3114 12005 3148
rect 11932 3080 11945 3114
rect 11979 3080 12005 3114
rect 11932 3046 12005 3080
rect 11932 3012 11945 3046
rect 11979 3012 12005 3046
rect 11932 2970 12005 3012
rect 12035 2991 12106 3170
rect 12136 3149 12189 3191
rect 12442 3178 12493 3190
rect 12442 3149 12450 3178
rect 12136 2991 12207 3149
rect 12035 2970 12088 2991
rect 12154 2949 12207 2991
rect 12237 3137 12297 3149
rect 12237 3103 12250 3137
rect 12284 3103 12297 3137
rect 12237 3069 12297 3103
rect 12237 3035 12250 3069
rect 12284 3035 12297 3069
rect 12237 3001 12297 3035
rect 12237 2967 12250 3001
rect 12284 2967 12297 3001
rect 12237 2949 12297 2967
rect 12327 3137 12394 3149
rect 12327 3103 12340 3137
rect 12374 3103 12394 3137
rect 12327 3045 12394 3103
rect 12327 3011 12340 3045
rect 12374 3011 12394 3045
rect 12327 2949 12394 3011
rect 12424 3144 12450 3149
rect 12484 3149 12493 3178
rect 13373 3182 13432 3194
rect 13062 3149 13181 3164
rect 12484 3144 12511 3149
rect 12424 2949 12511 3144
rect 12541 3110 12612 3149
rect 12541 3076 12554 3110
rect 12588 3076 12612 3110
rect 12541 2949 12612 3076
rect 12642 3113 12704 3149
rect 12642 3079 12655 3113
rect 12689 3079 12704 3113
rect 12642 2949 12704 3079
rect 12734 2949 12805 3149
rect 12835 3137 12895 3149
rect 12835 3103 12848 3137
rect 12882 3103 12895 3137
rect 12835 3026 12895 3103
rect 12835 2992 12848 3026
rect 12882 2992 12895 3026
rect 12835 2949 12895 2992
rect 12925 3137 13014 3149
rect 12925 3103 12967 3137
rect 13001 3103 13014 3137
rect 12925 3053 13014 3103
rect 12925 3019 12967 3053
rect 13001 3019 13014 3053
rect 12925 2949 13014 3019
rect 13044 3139 13181 3149
rect 13044 3105 13058 3139
rect 13092 3105 13133 3139
rect 13167 3105 13181 3139
rect 13044 2964 13181 3105
rect 13211 3152 13278 3164
rect 13211 3118 13232 3152
rect 13266 3118 13278 3152
rect 13211 3042 13278 3118
rect 13211 3008 13232 3042
rect 13266 3008 13278 3042
rect 13211 2964 13278 3008
rect 13373 3148 13385 3182
rect 13419 3148 13432 3182
rect 13373 3099 13432 3148
rect 13373 3065 13385 3099
rect 13419 3065 13432 3099
rect 13373 3016 13432 3065
rect 13373 2982 13385 3016
rect 13419 2982 13432 3016
rect 13373 2970 13432 2982
rect 13462 3182 13519 3194
rect 13462 3148 13475 3182
rect 13509 3148 13519 3182
rect 13462 3099 13519 3148
rect 13462 3065 13475 3099
rect 13509 3065 13519 3099
rect 13462 3016 13519 3065
rect 13462 2982 13475 3016
rect 13509 2982 13519 3016
rect 13462 2970 13519 2982
rect 13919 3180 13976 3192
rect 13919 3146 13929 3180
rect 13963 3146 13976 3180
rect 13919 3097 13976 3146
rect 13919 3063 13929 3097
rect 13963 3063 13976 3097
rect 13919 3014 13976 3063
rect 13919 2980 13929 3014
rect 13963 2980 13976 3014
rect 13044 2949 13097 2964
rect 13919 2968 13976 2980
rect 14006 3180 14061 3192
rect 14006 3146 14019 3180
rect 14053 3168 14061 3180
rect 14127 3168 14180 3189
rect 14053 3146 14079 3168
rect 14006 3112 14079 3146
rect 14006 3078 14019 3112
rect 14053 3078 14079 3112
rect 14006 3044 14079 3078
rect 14006 3010 14019 3044
rect 14053 3010 14079 3044
rect 14006 2968 14079 3010
rect 14109 2989 14180 3168
rect 14210 3147 14263 3189
rect 14516 3176 14567 3188
rect 14516 3147 14524 3176
rect 14210 2989 14281 3147
rect 14109 2968 14162 2989
rect 14228 2947 14281 2989
rect 14311 3135 14371 3147
rect 14311 3101 14324 3135
rect 14358 3101 14371 3135
rect 14311 3067 14371 3101
rect 14311 3033 14324 3067
rect 14358 3033 14371 3067
rect 14311 2999 14371 3033
rect 14311 2965 14324 2999
rect 14358 2965 14371 2999
rect 14311 2947 14371 2965
rect 14401 3135 14468 3147
rect 14401 3101 14414 3135
rect 14448 3101 14468 3135
rect 14401 3043 14468 3101
rect 14401 3009 14414 3043
rect 14448 3009 14468 3043
rect 14401 2947 14468 3009
rect 14498 3142 14524 3147
rect 14558 3147 14567 3176
rect 15447 3180 15506 3192
rect 15136 3147 15255 3162
rect 14558 3142 14585 3147
rect 14498 2947 14585 3142
rect 14615 3108 14686 3147
rect 14615 3074 14628 3108
rect 14662 3074 14686 3108
rect 14615 2947 14686 3074
rect 14716 3111 14778 3147
rect 14716 3077 14729 3111
rect 14763 3077 14778 3111
rect 14716 2947 14778 3077
rect 14808 2947 14879 3147
rect 14909 3135 14969 3147
rect 14909 3101 14922 3135
rect 14956 3101 14969 3135
rect 14909 3024 14969 3101
rect 14909 2990 14922 3024
rect 14956 2990 14969 3024
rect 14909 2947 14969 2990
rect 14999 3135 15088 3147
rect 14999 3101 15041 3135
rect 15075 3101 15088 3135
rect 14999 3051 15088 3101
rect 14999 3017 15041 3051
rect 15075 3017 15088 3051
rect 14999 2947 15088 3017
rect 15118 3137 15255 3147
rect 15118 3103 15132 3137
rect 15166 3103 15207 3137
rect 15241 3103 15255 3137
rect 15118 2962 15255 3103
rect 15285 3150 15352 3162
rect 15285 3116 15306 3150
rect 15340 3116 15352 3150
rect 15285 3040 15352 3116
rect 15285 3006 15306 3040
rect 15340 3006 15352 3040
rect 15285 2962 15352 3006
rect 15447 3146 15459 3180
rect 15493 3146 15506 3180
rect 15447 3097 15506 3146
rect 15447 3063 15459 3097
rect 15493 3063 15506 3097
rect 15447 3014 15506 3063
rect 15447 2980 15459 3014
rect 15493 2980 15506 3014
rect 15447 2968 15506 2980
rect 15536 3180 15593 3192
rect 15536 3146 15549 3180
rect 15583 3146 15593 3180
rect 15536 3097 15593 3146
rect 15536 3063 15549 3097
rect 15583 3063 15593 3097
rect 15536 3014 15593 3063
rect 15536 2980 15549 3014
rect 15583 2980 15593 3014
rect 15536 2968 15593 2980
rect 15981 3176 16038 3188
rect 15981 3142 15991 3176
rect 16025 3142 16038 3176
rect 15981 3093 16038 3142
rect 15981 3059 15991 3093
rect 16025 3059 16038 3093
rect 15981 3010 16038 3059
rect 15981 2976 15991 3010
rect 16025 2976 16038 3010
rect 15118 2947 15171 2962
rect 15981 2964 16038 2976
rect 16068 3176 16123 3188
rect 16068 3142 16081 3176
rect 16115 3164 16123 3176
rect 16189 3164 16242 3185
rect 16115 3142 16141 3164
rect 16068 3108 16141 3142
rect 16068 3074 16081 3108
rect 16115 3074 16141 3108
rect 16068 3040 16141 3074
rect 16068 3006 16081 3040
rect 16115 3006 16141 3040
rect 16068 2964 16141 3006
rect 16171 2985 16242 3164
rect 16272 3143 16325 3185
rect 16578 3172 16629 3184
rect 16578 3143 16586 3172
rect 16272 2985 16343 3143
rect 16171 2964 16224 2985
rect 16290 2943 16343 2985
rect 16373 3131 16433 3143
rect 16373 3097 16386 3131
rect 16420 3097 16433 3131
rect 16373 3063 16433 3097
rect 16373 3029 16386 3063
rect 16420 3029 16433 3063
rect 16373 2995 16433 3029
rect 16373 2961 16386 2995
rect 16420 2961 16433 2995
rect 16373 2943 16433 2961
rect 16463 3131 16530 3143
rect 16463 3097 16476 3131
rect 16510 3097 16530 3131
rect 16463 3039 16530 3097
rect 16463 3005 16476 3039
rect 16510 3005 16530 3039
rect 16463 2943 16530 3005
rect 16560 3138 16586 3143
rect 16620 3143 16629 3172
rect 17509 3176 17568 3188
rect 17198 3143 17317 3158
rect 16620 3138 16647 3143
rect 16560 2943 16647 3138
rect 16677 3104 16748 3143
rect 16677 3070 16690 3104
rect 16724 3070 16748 3104
rect 16677 2943 16748 3070
rect 16778 3107 16840 3143
rect 16778 3073 16791 3107
rect 16825 3073 16840 3107
rect 16778 2943 16840 3073
rect 16870 2943 16941 3143
rect 16971 3131 17031 3143
rect 16971 3097 16984 3131
rect 17018 3097 17031 3131
rect 16971 3020 17031 3097
rect 16971 2986 16984 3020
rect 17018 2986 17031 3020
rect 16971 2943 17031 2986
rect 17061 3131 17150 3143
rect 17061 3097 17103 3131
rect 17137 3097 17150 3131
rect 17061 3047 17150 3097
rect 17061 3013 17103 3047
rect 17137 3013 17150 3047
rect 17061 2943 17150 3013
rect 17180 3133 17317 3143
rect 17180 3099 17194 3133
rect 17228 3099 17269 3133
rect 17303 3099 17317 3133
rect 17180 2958 17317 3099
rect 17347 3146 17414 3158
rect 17347 3112 17368 3146
rect 17402 3112 17414 3146
rect 17347 3036 17414 3112
rect 17347 3002 17368 3036
rect 17402 3002 17414 3036
rect 17347 2958 17414 3002
rect 17509 3142 17521 3176
rect 17555 3142 17568 3176
rect 17509 3093 17568 3142
rect 17509 3059 17521 3093
rect 17555 3059 17568 3093
rect 17509 3010 17568 3059
rect 17509 2976 17521 3010
rect 17555 2976 17568 3010
rect 17509 2964 17568 2976
rect 17598 3176 17655 3188
rect 17598 3142 17611 3176
rect 17645 3142 17655 3176
rect 17598 3093 17655 3142
rect 17598 3059 17611 3093
rect 17645 3059 17655 3093
rect 17598 3010 17655 3059
rect 17598 2976 17611 3010
rect 17645 2976 17655 3010
rect 17598 2964 17655 2976
rect 17180 2943 17233 2958
<< ndiffc >>
rect 18198 5731 18232 5765
rect 18198 5663 18232 5697
rect 18282 5731 18316 5765
rect 18282 5663 18316 5697
rect 26340 5679 26374 5713
rect 26340 5611 26374 5645
rect 26424 5679 26458 5713
rect 26424 5611 26458 5645
rect 26508 5611 26542 5645
rect 26592 5679 26626 5713
rect 26592 5611 26626 5645
rect 26676 5611 26710 5645
rect 26760 5679 26794 5713
rect 26760 5611 26794 5645
rect 26844 5611 26878 5645
rect 26928 5679 26962 5713
rect 26928 5611 26962 5645
rect 27012 5611 27046 5645
rect 27096 5679 27130 5713
rect 27096 5611 27130 5645
rect 27180 5611 27214 5645
rect 27264 5679 27298 5713
rect 27264 5611 27298 5645
rect 27348 5611 27382 5645
rect 27432 5679 27466 5713
rect 27432 5611 27466 5645
rect 27516 5611 27550 5645
rect 27600 5679 27634 5713
rect 27600 5611 27634 5645
rect 27684 5679 27718 5713
rect 27684 5611 27718 5645
rect 28146 5661 28180 5695
rect 28146 5593 28180 5627
rect 28230 5661 28264 5695
rect 28230 5593 28264 5627
rect 28314 5593 28348 5627
rect 28398 5661 28432 5695
rect 28398 5593 28432 5627
rect 28482 5593 28516 5627
rect 28566 5661 28600 5695
rect 28566 5593 28600 5627
rect 28650 5593 28684 5627
rect 28734 5661 28768 5695
rect 28734 5593 28768 5627
rect 28818 5593 28852 5627
rect 28902 5661 28936 5695
rect 28902 5593 28936 5627
rect 28986 5593 29020 5627
rect 29070 5661 29104 5695
rect 29070 5593 29104 5627
rect 29154 5593 29188 5627
rect 29238 5661 29272 5695
rect 29238 5593 29272 5627
rect 29322 5593 29356 5627
rect 29406 5661 29440 5695
rect 29406 5593 29440 5627
rect 29490 5661 29524 5695
rect 29490 5593 29524 5627
rect 1537 2796 1571 2830
rect 1537 2706 1571 2740
rect 1641 2668 1675 2702
rect 1902 2713 1936 2747
rect 2018 2720 2052 2754
rect 2128 2668 2162 2702
rect 2230 2720 2264 2754
rect 2344 2712 2378 2746
rect 2523 2723 2557 2757
rect 2625 2671 2659 2705
rect 2719 2671 2753 2705
rect 2864 2664 2898 2698
rect 2966 2732 3000 2766
rect 3070 2724 3104 2758
rect 3156 2796 3190 2830
rect 3156 2706 3190 2740
rect 3599 2792 3633 2826
rect 3599 2702 3633 2736
rect 3703 2664 3737 2698
rect 3964 2709 3998 2743
rect 4080 2716 4114 2750
rect 4190 2664 4224 2698
rect 4292 2716 4326 2750
rect 4406 2708 4440 2742
rect 4585 2719 4619 2753
rect 4687 2667 4721 2701
rect 4781 2667 4815 2701
rect 4926 2660 4960 2694
rect 5028 2728 5062 2762
rect 5132 2720 5166 2754
rect 5218 2792 5252 2826
rect 5218 2702 5252 2736
rect 5673 2790 5707 2824
rect 5673 2700 5707 2734
rect 5777 2662 5811 2696
rect 6038 2707 6072 2741
rect 6154 2714 6188 2748
rect 6264 2662 6298 2696
rect 6366 2714 6400 2748
rect 6480 2706 6514 2740
rect 6659 2717 6693 2751
rect 6761 2665 6795 2699
rect 6855 2665 6889 2699
rect 7000 2658 7034 2692
rect 7102 2726 7136 2760
rect 7206 2718 7240 2752
rect 7292 2790 7326 2824
rect 7292 2700 7326 2734
rect 7735 2786 7769 2820
rect 7735 2696 7769 2730
rect 7839 2658 7873 2692
rect 8100 2703 8134 2737
rect 8216 2710 8250 2744
rect 8326 2658 8360 2692
rect 8428 2710 8462 2744
rect 8542 2702 8576 2736
rect 8721 2713 8755 2747
rect 8823 2661 8857 2695
rect 8917 2661 8951 2695
rect 9062 2654 9096 2688
rect 9164 2722 9198 2756
rect 9268 2714 9302 2748
rect 9354 2786 9388 2820
rect 9354 2696 9388 2730
rect 9795 2782 9829 2816
rect 9795 2692 9829 2726
rect 9899 2654 9933 2688
rect 10160 2699 10194 2733
rect 10276 2706 10310 2740
rect 10386 2654 10420 2688
rect 10488 2706 10522 2740
rect 10602 2698 10636 2732
rect 10781 2709 10815 2743
rect 10883 2657 10917 2691
rect 10977 2657 11011 2691
rect 11122 2650 11156 2684
rect 11224 2718 11258 2752
rect 11328 2710 11362 2744
rect 11414 2782 11448 2816
rect 11414 2692 11448 2726
rect 11857 2778 11891 2812
rect 11857 2688 11891 2722
rect 11961 2650 11995 2684
rect 12222 2695 12256 2729
rect 12338 2702 12372 2736
rect 12448 2650 12482 2684
rect 12550 2702 12584 2736
rect 12664 2694 12698 2728
rect 12843 2705 12877 2739
rect 12945 2653 12979 2687
rect 13039 2653 13073 2687
rect 13184 2646 13218 2680
rect 13286 2714 13320 2748
rect 13390 2706 13424 2740
rect 13476 2778 13510 2812
rect 13476 2688 13510 2722
rect 13931 2776 13965 2810
rect 13931 2686 13965 2720
rect 14035 2648 14069 2682
rect 14296 2693 14330 2727
rect 14412 2700 14446 2734
rect 14522 2648 14556 2682
rect 14624 2700 14658 2734
rect 14738 2692 14772 2726
rect 14917 2703 14951 2737
rect 15019 2651 15053 2685
rect 15113 2651 15147 2685
rect 15258 2644 15292 2678
rect 15360 2712 15394 2746
rect 15464 2704 15498 2738
rect 15550 2776 15584 2810
rect 15550 2686 15584 2720
rect 15993 2772 16027 2806
rect 15993 2682 16027 2716
rect 16097 2644 16131 2678
rect 16358 2689 16392 2723
rect 16474 2696 16508 2730
rect 16584 2644 16618 2678
rect 16686 2696 16720 2730
rect 16800 2688 16834 2722
rect 16979 2699 17013 2733
rect 17081 2647 17115 2681
rect 17175 2647 17209 2681
rect 17320 2640 17354 2674
rect 17422 2708 17456 2742
rect 17526 2700 17560 2734
rect 17612 2772 17646 2806
rect 17612 2682 17646 2716
<< pdiffc >>
rect 18198 6051 18232 6085
rect 18198 5983 18232 6017
rect 18198 5915 18232 5949
rect 18282 6051 18316 6085
rect 18282 5983 18316 6017
rect 18282 5915 18316 5949
rect 26340 6003 26374 6037
rect 26340 5935 26374 5969
rect 26340 5865 26374 5899
rect 26424 6003 26458 6037
rect 26424 5935 26458 5969
rect 26424 5865 26458 5899
rect 26508 6003 26542 6037
rect 26508 5935 26542 5969
rect 26592 6003 26626 6037
rect 26592 5935 26626 5969
rect 26592 5865 26626 5899
rect 26676 6003 26710 6037
rect 26676 5935 26710 5969
rect 26760 6003 26794 6037
rect 26760 5935 26794 5969
rect 26760 5865 26794 5899
rect 26844 6003 26878 6037
rect 26844 5935 26878 5969
rect 26928 6003 26962 6037
rect 26928 5935 26962 5969
rect 26928 5865 26962 5899
rect 27012 6003 27046 6037
rect 27012 5935 27046 5969
rect 27096 6003 27130 6037
rect 27096 5935 27130 5969
rect 27096 5865 27130 5899
rect 27180 6003 27214 6037
rect 27180 5935 27214 5969
rect 27264 6003 27298 6037
rect 27264 5935 27298 5969
rect 27264 5865 27298 5899
rect 27348 6003 27382 6037
rect 27348 5935 27382 5969
rect 27432 6003 27466 6037
rect 27432 5935 27466 5969
rect 27432 5865 27466 5899
rect 27516 6003 27550 6037
rect 27516 5935 27550 5969
rect 27600 6003 27634 6037
rect 27600 5935 27634 5969
rect 27600 5865 27634 5899
rect 27684 6003 27718 6037
rect 27684 5935 27718 5969
rect 28146 5985 28180 6019
rect 28146 5917 28180 5951
rect 28146 5847 28180 5881
rect 28230 5985 28264 6019
rect 28230 5917 28264 5951
rect 28230 5847 28264 5881
rect 28314 5985 28348 6019
rect 28314 5917 28348 5951
rect 28398 5985 28432 6019
rect 28398 5917 28432 5951
rect 28398 5847 28432 5881
rect 28482 5985 28516 6019
rect 28482 5917 28516 5951
rect 28566 5985 28600 6019
rect 28566 5917 28600 5951
rect 28566 5847 28600 5881
rect 28650 5985 28684 6019
rect 28650 5917 28684 5951
rect 28734 5985 28768 6019
rect 28734 5917 28768 5951
rect 28734 5847 28768 5881
rect 28818 5985 28852 6019
rect 28818 5917 28852 5951
rect 28902 5985 28936 6019
rect 28902 5917 28936 5951
rect 28902 5847 28936 5881
rect 28986 5985 29020 6019
rect 28986 5917 29020 5951
rect 29070 5985 29104 6019
rect 29070 5917 29104 5951
rect 29070 5847 29104 5881
rect 29154 5985 29188 6019
rect 29154 5917 29188 5951
rect 29238 5985 29272 6019
rect 29238 5917 29272 5951
rect 29238 5847 29272 5881
rect 29322 5985 29356 6019
rect 29322 5917 29356 5951
rect 29406 5985 29440 6019
rect 29406 5917 29440 5951
rect 29406 5847 29440 5881
rect 29490 5985 29524 6019
rect 29490 5917 29524 5951
rect 1535 3166 1569 3200
rect 1535 3083 1569 3117
rect 1535 3000 1569 3034
rect 1625 3166 1659 3200
rect 1625 3098 1659 3132
rect 1625 3030 1659 3064
rect 1930 3121 1964 3155
rect 1930 3053 1964 3087
rect 1930 2985 1964 3019
rect 2020 3121 2054 3155
rect 2020 3029 2054 3063
rect 2130 3162 2164 3196
rect 2234 3094 2268 3128
rect 2335 3097 2369 3131
rect 2528 3121 2562 3155
rect 2528 3010 2562 3044
rect 2647 3121 2681 3155
rect 2647 3037 2681 3071
rect 2738 3123 2772 3157
rect 2813 3123 2847 3157
rect 2912 3136 2946 3170
rect 2912 3026 2946 3060
rect 3065 3166 3099 3200
rect 3065 3083 3099 3117
rect 3065 3000 3099 3034
rect 3155 3166 3189 3200
rect 3155 3083 3189 3117
rect 3155 3000 3189 3034
rect 3597 3162 3631 3196
rect 3597 3079 3631 3113
rect 3597 2996 3631 3030
rect 3687 3162 3721 3196
rect 3687 3094 3721 3128
rect 3687 3026 3721 3060
rect 3992 3117 4026 3151
rect 3992 3049 4026 3083
rect 3992 2981 4026 3015
rect 4082 3117 4116 3151
rect 4082 3025 4116 3059
rect 4192 3158 4226 3192
rect 4296 3090 4330 3124
rect 4397 3093 4431 3127
rect 4590 3117 4624 3151
rect 4590 3006 4624 3040
rect 4709 3117 4743 3151
rect 4709 3033 4743 3067
rect 4800 3119 4834 3153
rect 4875 3119 4909 3153
rect 4974 3132 5008 3166
rect 4974 3022 5008 3056
rect 5127 3162 5161 3196
rect 5127 3079 5161 3113
rect 5127 2996 5161 3030
rect 5217 3162 5251 3196
rect 5217 3079 5251 3113
rect 5217 2996 5251 3030
rect 5671 3160 5705 3194
rect 5671 3077 5705 3111
rect 5671 2994 5705 3028
rect 5761 3160 5795 3194
rect 5761 3092 5795 3126
rect 5761 3024 5795 3058
rect 6066 3115 6100 3149
rect 6066 3047 6100 3081
rect 6066 2979 6100 3013
rect 6156 3115 6190 3149
rect 6156 3023 6190 3057
rect 6266 3156 6300 3190
rect 6370 3088 6404 3122
rect 6471 3091 6505 3125
rect 6664 3115 6698 3149
rect 6664 3004 6698 3038
rect 6783 3115 6817 3149
rect 6783 3031 6817 3065
rect 6874 3117 6908 3151
rect 6949 3117 6983 3151
rect 7048 3130 7082 3164
rect 7048 3020 7082 3054
rect 7201 3160 7235 3194
rect 7201 3077 7235 3111
rect 7201 2994 7235 3028
rect 7291 3160 7325 3194
rect 7291 3077 7325 3111
rect 7291 2994 7325 3028
rect 7733 3156 7767 3190
rect 7733 3073 7767 3107
rect 7733 2990 7767 3024
rect 7823 3156 7857 3190
rect 7823 3088 7857 3122
rect 7823 3020 7857 3054
rect 8128 3111 8162 3145
rect 8128 3043 8162 3077
rect 8128 2975 8162 3009
rect 8218 3111 8252 3145
rect 8218 3019 8252 3053
rect 8328 3152 8362 3186
rect 8432 3084 8466 3118
rect 8533 3087 8567 3121
rect 8726 3111 8760 3145
rect 8726 3000 8760 3034
rect 8845 3111 8879 3145
rect 8845 3027 8879 3061
rect 8936 3113 8970 3147
rect 9011 3113 9045 3147
rect 9110 3126 9144 3160
rect 9110 3016 9144 3050
rect 9263 3156 9297 3190
rect 9263 3073 9297 3107
rect 9263 2990 9297 3024
rect 9353 3156 9387 3190
rect 9353 3073 9387 3107
rect 9353 2990 9387 3024
rect 9793 3152 9827 3186
rect 9793 3069 9827 3103
rect 9793 2986 9827 3020
rect 9883 3152 9917 3186
rect 9883 3084 9917 3118
rect 9883 3016 9917 3050
rect 10188 3107 10222 3141
rect 10188 3039 10222 3073
rect 10188 2971 10222 3005
rect 10278 3107 10312 3141
rect 10278 3015 10312 3049
rect 10388 3148 10422 3182
rect 10492 3080 10526 3114
rect 10593 3083 10627 3117
rect 10786 3107 10820 3141
rect 10786 2996 10820 3030
rect 10905 3107 10939 3141
rect 10905 3023 10939 3057
rect 10996 3109 11030 3143
rect 11071 3109 11105 3143
rect 11170 3122 11204 3156
rect 11170 3012 11204 3046
rect 11323 3152 11357 3186
rect 11323 3069 11357 3103
rect 11323 2986 11357 3020
rect 11413 3152 11447 3186
rect 11413 3069 11447 3103
rect 11413 2986 11447 3020
rect 11855 3148 11889 3182
rect 11855 3065 11889 3099
rect 11855 2982 11889 3016
rect 11945 3148 11979 3182
rect 11945 3080 11979 3114
rect 11945 3012 11979 3046
rect 12250 3103 12284 3137
rect 12250 3035 12284 3069
rect 12250 2967 12284 3001
rect 12340 3103 12374 3137
rect 12340 3011 12374 3045
rect 12450 3144 12484 3178
rect 12554 3076 12588 3110
rect 12655 3079 12689 3113
rect 12848 3103 12882 3137
rect 12848 2992 12882 3026
rect 12967 3103 13001 3137
rect 12967 3019 13001 3053
rect 13058 3105 13092 3139
rect 13133 3105 13167 3139
rect 13232 3118 13266 3152
rect 13232 3008 13266 3042
rect 13385 3148 13419 3182
rect 13385 3065 13419 3099
rect 13385 2982 13419 3016
rect 13475 3148 13509 3182
rect 13475 3065 13509 3099
rect 13475 2982 13509 3016
rect 13929 3146 13963 3180
rect 13929 3063 13963 3097
rect 13929 2980 13963 3014
rect 14019 3146 14053 3180
rect 14019 3078 14053 3112
rect 14019 3010 14053 3044
rect 14324 3101 14358 3135
rect 14324 3033 14358 3067
rect 14324 2965 14358 2999
rect 14414 3101 14448 3135
rect 14414 3009 14448 3043
rect 14524 3142 14558 3176
rect 14628 3074 14662 3108
rect 14729 3077 14763 3111
rect 14922 3101 14956 3135
rect 14922 2990 14956 3024
rect 15041 3101 15075 3135
rect 15041 3017 15075 3051
rect 15132 3103 15166 3137
rect 15207 3103 15241 3137
rect 15306 3116 15340 3150
rect 15306 3006 15340 3040
rect 15459 3146 15493 3180
rect 15459 3063 15493 3097
rect 15459 2980 15493 3014
rect 15549 3146 15583 3180
rect 15549 3063 15583 3097
rect 15549 2980 15583 3014
rect 15991 3142 16025 3176
rect 15991 3059 16025 3093
rect 15991 2976 16025 3010
rect 16081 3142 16115 3176
rect 16081 3074 16115 3108
rect 16081 3006 16115 3040
rect 16386 3097 16420 3131
rect 16386 3029 16420 3063
rect 16386 2961 16420 2995
rect 16476 3097 16510 3131
rect 16476 3005 16510 3039
rect 16586 3138 16620 3172
rect 16690 3070 16724 3104
rect 16791 3073 16825 3107
rect 16984 3097 17018 3131
rect 16984 2986 17018 3020
rect 17103 3097 17137 3131
rect 17103 3013 17137 3047
rect 17194 3099 17228 3133
rect 17269 3099 17303 3133
rect 17368 3112 17402 3146
rect 17368 3002 17402 3036
rect 17521 3142 17555 3176
rect 17521 3059 17555 3093
rect 17521 2976 17555 3010
rect 17611 3142 17645 3176
rect 17611 3059 17645 3093
rect 17611 2976 17645 3010
<< poly >>
rect 18242 6097 18272 6123
rect 26384 6049 26414 6075
rect 26468 6049 26498 6075
rect 26552 6049 26582 6075
rect 26636 6049 26666 6075
rect 26720 6049 26750 6075
rect 26804 6049 26834 6075
rect 26888 6049 26918 6075
rect 26972 6049 27002 6075
rect 27056 6049 27086 6075
rect 27140 6049 27170 6075
rect 27224 6049 27254 6075
rect 27308 6049 27338 6075
rect 27392 6049 27422 6075
rect 27476 6049 27506 6075
rect 27560 6049 27590 6075
rect 27644 6049 27674 6075
rect 18242 5865 18272 5897
rect 18186 5849 18272 5865
rect 28190 6031 28220 6057
rect 28274 6031 28304 6057
rect 28358 6031 28388 6057
rect 28442 6031 28472 6057
rect 28526 6031 28556 6057
rect 28610 6031 28640 6057
rect 28694 6031 28724 6057
rect 28778 6031 28808 6057
rect 28862 6031 28892 6057
rect 28946 6031 28976 6057
rect 29030 6031 29060 6057
rect 29114 6031 29144 6057
rect 29198 6031 29228 6057
rect 29282 6031 29312 6057
rect 29366 6031 29396 6057
rect 29450 6031 29480 6057
rect 18186 5815 18202 5849
rect 18236 5815 18272 5849
rect 26384 5817 26414 5849
rect 26468 5817 26498 5849
rect 26552 5817 26582 5849
rect 26636 5817 26666 5849
rect 26720 5817 26750 5849
rect 26804 5817 26834 5849
rect 26888 5817 26918 5849
rect 26972 5817 27002 5849
rect 27056 5817 27086 5849
rect 27140 5817 27170 5849
rect 27224 5817 27254 5849
rect 27308 5817 27338 5849
rect 27392 5817 27422 5849
rect 27476 5817 27506 5849
rect 27560 5817 27590 5849
rect 27644 5817 27674 5849
rect 18186 5799 18272 5815
rect 18242 5777 18272 5799
rect 26318 5801 27674 5817
rect 26318 5767 26334 5801
rect 26368 5767 26508 5801
rect 26542 5767 26676 5801
rect 26710 5767 26845 5801
rect 26879 5767 27012 5801
rect 27046 5767 27180 5801
rect 27214 5767 27347 5801
rect 27381 5767 27674 5801
rect 28190 5799 28220 5831
rect 28274 5799 28304 5831
rect 28358 5799 28388 5831
rect 28442 5799 28472 5831
rect 28526 5799 28556 5831
rect 28610 5799 28640 5831
rect 28694 5799 28724 5831
rect 28778 5799 28808 5831
rect 28862 5799 28892 5831
rect 28946 5799 28976 5831
rect 29030 5799 29060 5831
rect 29114 5799 29144 5831
rect 29198 5799 29228 5831
rect 29282 5799 29312 5831
rect 29366 5799 29396 5831
rect 29450 5799 29480 5831
rect 26318 5751 27674 5767
rect 26384 5729 26414 5751
rect 26468 5729 26498 5751
rect 26552 5729 26582 5751
rect 26636 5729 26666 5751
rect 26720 5729 26750 5751
rect 26804 5729 26834 5751
rect 26888 5729 26918 5751
rect 26972 5729 27002 5751
rect 27056 5729 27086 5751
rect 27140 5729 27170 5751
rect 27224 5729 27254 5751
rect 27308 5729 27338 5751
rect 27392 5729 27422 5751
rect 27476 5729 27506 5751
rect 27560 5729 27590 5751
rect 27644 5729 27674 5751
rect 28124 5783 29480 5799
rect 28124 5749 28140 5783
rect 28174 5749 28314 5783
rect 28348 5749 28482 5783
rect 28516 5749 28651 5783
rect 28685 5749 28818 5783
rect 28852 5749 28986 5783
rect 29020 5749 29153 5783
rect 29187 5749 29480 5783
rect 28124 5733 29480 5749
rect 18242 5621 18272 5647
rect 28190 5711 28220 5733
rect 28274 5711 28304 5733
rect 28358 5711 28388 5733
rect 28442 5711 28472 5733
rect 28526 5711 28556 5733
rect 28610 5711 28640 5733
rect 28694 5711 28724 5733
rect 28778 5711 28808 5733
rect 28862 5711 28892 5733
rect 28946 5711 28976 5733
rect 29030 5711 29060 5733
rect 29114 5711 29144 5733
rect 29198 5711 29228 5733
rect 29282 5711 29312 5733
rect 29366 5711 29396 5733
rect 29450 5711 29480 5733
rect 26384 5573 26414 5599
rect 26468 5573 26498 5599
rect 26552 5573 26582 5599
rect 26636 5573 26666 5599
rect 26720 5573 26750 5599
rect 26804 5573 26834 5599
rect 26888 5573 26918 5599
rect 26972 5573 27002 5599
rect 27056 5573 27086 5599
rect 27140 5573 27170 5599
rect 27224 5573 27254 5599
rect 27308 5573 27338 5599
rect 27392 5573 27422 5599
rect 27476 5573 27506 5599
rect 27560 5573 27590 5599
rect 27644 5573 27674 5599
rect 28190 5555 28220 5581
rect 28274 5555 28304 5581
rect 28358 5555 28388 5581
rect 28442 5555 28472 5581
rect 28526 5555 28556 5581
rect 28610 5555 28640 5581
rect 28694 5555 28724 5581
rect 28778 5555 28808 5581
rect 28862 5555 28892 5581
rect 28946 5555 28976 5581
rect 29030 5555 29060 5581
rect 29114 5555 29144 5581
rect 29198 5555 29228 5581
rect 29282 5555 29312 5581
rect 29366 5555 29396 5581
rect 29450 5555 29480 5581
rect 1582 3212 1612 3238
rect 1783 3235 2894 3265
rect 1783 3224 1819 3235
rect 1685 3188 1715 3214
rect 1786 3209 1816 3224
rect 1887 3167 1917 3193
rect 1977 3167 2007 3193
rect 2071 3182 2107 3235
rect 2074 3167 2104 3182
rect 1786 2994 1816 3009
rect 1582 2973 1612 2988
rect 1685 2973 1715 2988
rect 1579 2946 1615 2973
rect 1567 2930 1633 2946
rect 1682 2930 1718 2973
rect 1783 2963 1819 2994
rect 2191 3167 2221 3193
rect 2292 3167 2322 3193
rect 2384 3167 2414 3193
rect 2482 3182 2518 3235
rect 2858 3197 2894 3235
rect 3112 3212 3142 3238
rect 2485 3167 2515 3182
rect 2575 3167 2605 3193
rect 2694 3167 2724 3193
rect 2861 3182 2891 3197
rect 3644 3208 3674 3234
rect 3845 3231 4956 3261
rect 3845 3220 3881 3231
rect 2861 2967 2891 2982
rect 3112 2973 3142 2988
rect 3747 3184 3777 3210
rect 3848 3205 3878 3220
rect 3949 3163 3979 3189
rect 4039 3163 4069 3189
rect 4133 3178 4169 3231
rect 4136 3163 4166 3178
rect 3848 2990 3878 3005
rect 1567 2896 1583 2930
rect 1617 2896 1633 2930
rect 1567 2880 1633 2896
rect 1675 2914 1741 2930
rect 1675 2880 1691 2914
rect 1725 2880 1741 2914
rect 1582 2842 1612 2880
rect 1675 2864 1741 2880
rect 1705 2823 1735 2864
rect 1783 2823 1813 2963
rect 1887 2952 1917 2967
rect 1977 2952 2007 2967
rect 2074 2952 2104 2967
rect 2191 2952 2221 2967
rect 2292 2952 2322 2967
rect 2384 2952 2414 2967
rect 2485 2952 2515 2967
rect 2575 2952 2605 2967
rect 2694 2952 2724 2967
rect 1884 2935 1920 2952
rect 1974 2935 2010 2952
rect 1855 2919 1921 2935
rect 1855 2885 1871 2919
rect 1905 2885 1921 2919
rect 1855 2869 1921 2885
rect 1963 2919 2029 2935
rect 1963 2885 1979 2919
rect 2013 2885 2029 2919
rect 1963 2869 2029 2885
rect 1861 2823 1891 2869
rect 1969 2823 1999 2869
rect 2071 2838 2107 2952
rect 2188 2911 2224 2952
rect 2289 2935 2325 2952
rect 2158 2895 2224 2911
rect 2158 2861 2174 2895
rect 2208 2861 2224 2895
rect 2266 2919 2332 2935
rect 2266 2885 2282 2919
rect 2316 2885 2332 2919
rect 2381 2911 2417 2952
rect 2266 2869 2332 2885
rect 2374 2895 2440 2911
rect 2158 2845 2224 2861
rect 2071 2823 2101 2838
rect 2189 2823 2219 2845
rect 2275 2823 2305 2869
rect 2374 2861 2390 2895
rect 2424 2861 2440 2895
rect 2374 2845 2440 2861
rect 2404 2823 2434 2845
rect 2482 2838 2518 2952
rect 2572 2935 2608 2952
rect 2691 2935 2727 2952
rect 2858 2950 2894 2967
rect 2560 2919 2626 2935
rect 2560 2885 2576 2919
rect 2610 2885 2626 2919
rect 2560 2869 2626 2885
rect 2674 2919 2740 2935
rect 2674 2885 2690 2919
rect 2724 2885 2740 2919
rect 2674 2872 2740 2885
rect 2858 2934 2992 2950
rect 2858 2900 2874 2934
rect 2908 2900 2942 2934
rect 2976 2900 2992 2934
rect 3109 2930 3145 2973
rect 3644 2969 3674 2984
rect 3747 2969 3777 2984
rect 3641 2942 3677 2969
rect 2858 2884 2992 2900
rect 3040 2914 3145 2930
rect 2482 2823 2512 2838
rect 2568 2823 2598 2869
rect 2674 2842 2810 2872
rect 2780 2823 2810 2842
rect 2925 2823 2955 2884
rect 3040 2880 3056 2914
rect 3090 2880 3145 2914
rect 3040 2864 3145 2880
rect 3629 2926 3695 2942
rect 3744 2926 3780 2969
rect 3845 2959 3881 2990
rect 4253 3163 4283 3189
rect 4354 3163 4384 3189
rect 4446 3163 4476 3189
rect 4544 3178 4580 3231
rect 4920 3193 4956 3231
rect 5174 3208 5204 3234
rect 4547 3163 4577 3178
rect 4637 3163 4667 3189
rect 4756 3163 4786 3189
rect 4923 3178 4953 3193
rect 5718 3206 5748 3232
rect 5919 3229 7030 3259
rect 5919 3218 5955 3229
rect 4923 2963 4953 2978
rect 5174 2969 5204 2984
rect 5821 3182 5851 3208
rect 5922 3203 5952 3218
rect 6023 3161 6053 3187
rect 6113 3161 6143 3187
rect 6207 3176 6243 3229
rect 6210 3161 6240 3176
rect 5922 2988 5952 3003
rect 3629 2892 3645 2926
rect 3679 2892 3695 2926
rect 3629 2876 3695 2892
rect 3737 2910 3803 2926
rect 3737 2876 3753 2910
rect 3787 2876 3803 2910
rect 3115 2842 3145 2864
rect 1582 2668 1612 2694
rect 1705 2669 1735 2695
rect 1783 2669 1813 2695
rect 1861 2669 1891 2695
rect 1969 2669 1999 2695
rect 2071 2669 2101 2695
rect 2189 2669 2219 2695
rect 2275 2669 2305 2695
rect 2404 2669 2434 2695
rect 2482 2669 2512 2695
rect 2568 2669 2598 2695
rect 2780 2669 2810 2695
rect 2925 2669 2955 2695
rect 3644 2838 3674 2876
rect 3737 2860 3803 2876
rect 3115 2668 3145 2694
rect 3767 2819 3797 2860
rect 3845 2819 3875 2959
rect 3949 2948 3979 2963
rect 4039 2948 4069 2963
rect 4136 2948 4166 2963
rect 4253 2948 4283 2963
rect 4354 2948 4384 2963
rect 4446 2948 4476 2963
rect 4547 2948 4577 2963
rect 4637 2948 4667 2963
rect 4756 2948 4786 2963
rect 3946 2931 3982 2948
rect 4036 2931 4072 2948
rect 3917 2915 3983 2931
rect 3917 2881 3933 2915
rect 3967 2881 3983 2915
rect 3917 2865 3983 2881
rect 4025 2915 4091 2931
rect 4025 2881 4041 2915
rect 4075 2881 4091 2915
rect 4025 2865 4091 2881
rect 3923 2819 3953 2865
rect 4031 2819 4061 2865
rect 4133 2834 4169 2948
rect 4250 2907 4286 2948
rect 4351 2931 4387 2948
rect 4220 2891 4286 2907
rect 4220 2857 4236 2891
rect 4270 2857 4286 2891
rect 4328 2915 4394 2931
rect 4328 2881 4344 2915
rect 4378 2881 4394 2915
rect 4443 2907 4479 2948
rect 4328 2865 4394 2881
rect 4436 2891 4502 2907
rect 4220 2841 4286 2857
rect 4133 2819 4163 2834
rect 4251 2819 4281 2841
rect 4337 2819 4367 2865
rect 4436 2857 4452 2891
rect 4486 2857 4502 2891
rect 4436 2841 4502 2857
rect 4466 2819 4496 2841
rect 4544 2834 4580 2948
rect 4634 2931 4670 2948
rect 4753 2931 4789 2948
rect 4920 2946 4956 2963
rect 4622 2915 4688 2931
rect 4622 2881 4638 2915
rect 4672 2881 4688 2915
rect 4622 2865 4688 2881
rect 4736 2915 4802 2931
rect 4736 2881 4752 2915
rect 4786 2881 4802 2915
rect 4736 2868 4802 2881
rect 4920 2930 5054 2946
rect 4920 2896 4936 2930
rect 4970 2896 5004 2930
rect 5038 2896 5054 2930
rect 5171 2926 5207 2969
rect 5718 2967 5748 2982
rect 5821 2967 5851 2982
rect 5715 2940 5751 2967
rect 4920 2880 5054 2896
rect 5102 2910 5207 2926
rect 4544 2819 4574 2834
rect 4630 2819 4660 2865
rect 4736 2838 4872 2868
rect 4842 2819 4872 2838
rect 4987 2819 5017 2880
rect 5102 2876 5118 2910
rect 5152 2876 5207 2910
rect 5102 2860 5207 2876
rect 5703 2924 5769 2940
rect 5818 2924 5854 2967
rect 5919 2957 5955 2988
rect 6327 3161 6357 3187
rect 6428 3161 6458 3187
rect 6520 3161 6550 3187
rect 6618 3176 6654 3229
rect 6994 3191 7030 3229
rect 7248 3206 7278 3232
rect 6621 3161 6651 3176
rect 6711 3161 6741 3187
rect 6830 3161 6860 3187
rect 6997 3176 7027 3191
rect 7780 3202 7810 3228
rect 7981 3225 9092 3255
rect 7981 3214 8017 3225
rect 6997 2961 7027 2976
rect 7248 2967 7278 2982
rect 7883 3178 7913 3204
rect 7984 3199 8014 3214
rect 8085 3157 8115 3183
rect 8175 3157 8205 3183
rect 8269 3172 8305 3225
rect 8272 3157 8302 3172
rect 7984 2984 8014 2999
rect 5703 2890 5719 2924
rect 5753 2890 5769 2924
rect 5703 2874 5769 2890
rect 5811 2908 5877 2924
rect 5811 2874 5827 2908
rect 5861 2874 5877 2908
rect 5177 2838 5207 2860
rect 3644 2664 3674 2690
rect 3767 2665 3797 2691
rect 3845 2665 3875 2691
rect 3923 2665 3953 2691
rect 4031 2665 4061 2691
rect 4133 2665 4163 2691
rect 4251 2665 4281 2691
rect 4337 2665 4367 2691
rect 4466 2665 4496 2691
rect 4544 2665 4574 2691
rect 4630 2665 4660 2691
rect 4842 2665 4872 2691
rect 4987 2665 5017 2691
rect 5718 2836 5748 2874
rect 5811 2858 5877 2874
rect 5177 2664 5207 2690
rect 5841 2817 5871 2858
rect 5919 2817 5949 2957
rect 6023 2946 6053 2961
rect 6113 2946 6143 2961
rect 6210 2946 6240 2961
rect 6327 2946 6357 2961
rect 6428 2946 6458 2961
rect 6520 2946 6550 2961
rect 6621 2946 6651 2961
rect 6711 2946 6741 2961
rect 6830 2946 6860 2961
rect 6020 2929 6056 2946
rect 6110 2929 6146 2946
rect 5991 2913 6057 2929
rect 5991 2879 6007 2913
rect 6041 2879 6057 2913
rect 5991 2863 6057 2879
rect 6099 2913 6165 2929
rect 6099 2879 6115 2913
rect 6149 2879 6165 2913
rect 6099 2863 6165 2879
rect 5997 2817 6027 2863
rect 6105 2817 6135 2863
rect 6207 2832 6243 2946
rect 6324 2905 6360 2946
rect 6425 2929 6461 2946
rect 6294 2889 6360 2905
rect 6294 2855 6310 2889
rect 6344 2855 6360 2889
rect 6402 2913 6468 2929
rect 6402 2879 6418 2913
rect 6452 2879 6468 2913
rect 6517 2905 6553 2946
rect 6402 2863 6468 2879
rect 6510 2889 6576 2905
rect 6294 2839 6360 2855
rect 6207 2817 6237 2832
rect 6325 2817 6355 2839
rect 6411 2817 6441 2863
rect 6510 2855 6526 2889
rect 6560 2855 6576 2889
rect 6510 2839 6576 2855
rect 6540 2817 6570 2839
rect 6618 2832 6654 2946
rect 6708 2929 6744 2946
rect 6827 2929 6863 2946
rect 6994 2944 7030 2961
rect 6696 2913 6762 2929
rect 6696 2879 6712 2913
rect 6746 2879 6762 2913
rect 6696 2863 6762 2879
rect 6810 2913 6876 2929
rect 6810 2879 6826 2913
rect 6860 2879 6876 2913
rect 6810 2866 6876 2879
rect 6994 2928 7128 2944
rect 6994 2894 7010 2928
rect 7044 2894 7078 2928
rect 7112 2894 7128 2928
rect 7245 2924 7281 2967
rect 7780 2963 7810 2978
rect 7883 2963 7913 2978
rect 7777 2936 7813 2963
rect 6994 2878 7128 2894
rect 7176 2908 7281 2924
rect 6618 2817 6648 2832
rect 6704 2817 6734 2863
rect 6810 2836 6946 2866
rect 6916 2817 6946 2836
rect 7061 2817 7091 2878
rect 7176 2874 7192 2908
rect 7226 2874 7281 2908
rect 7176 2858 7281 2874
rect 7765 2920 7831 2936
rect 7880 2920 7916 2963
rect 7981 2953 8017 2984
rect 8389 3157 8419 3183
rect 8490 3157 8520 3183
rect 8582 3157 8612 3183
rect 8680 3172 8716 3225
rect 9056 3187 9092 3225
rect 9310 3202 9340 3228
rect 8683 3157 8713 3172
rect 8773 3157 8803 3183
rect 8892 3157 8922 3183
rect 9059 3172 9089 3187
rect 9840 3198 9870 3224
rect 10041 3221 11152 3251
rect 10041 3210 10077 3221
rect 9059 2957 9089 2972
rect 9310 2963 9340 2978
rect 9943 3174 9973 3200
rect 10044 3195 10074 3210
rect 10145 3153 10175 3179
rect 10235 3153 10265 3179
rect 10329 3168 10365 3221
rect 10332 3153 10362 3168
rect 10044 2980 10074 2995
rect 7765 2886 7781 2920
rect 7815 2886 7831 2920
rect 7765 2870 7831 2886
rect 7873 2904 7939 2920
rect 7873 2870 7889 2904
rect 7923 2870 7939 2904
rect 7251 2836 7281 2858
rect 5718 2662 5748 2688
rect 5841 2663 5871 2689
rect 5919 2663 5949 2689
rect 5997 2663 6027 2689
rect 6105 2663 6135 2689
rect 6207 2663 6237 2689
rect 6325 2663 6355 2689
rect 6411 2663 6441 2689
rect 6540 2663 6570 2689
rect 6618 2663 6648 2689
rect 6704 2663 6734 2689
rect 6916 2663 6946 2689
rect 7061 2663 7091 2689
rect 7780 2832 7810 2870
rect 7873 2854 7939 2870
rect 7251 2662 7281 2688
rect 7903 2813 7933 2854
rect 7981 2813 8011 2953
rect 8085 2942 8115 2957
rect 8175 2942 8205 2957
rect 8272 2942 8302 2957
rect 8389 2942 8419 2957
rect 8490 2942 8520 2957
rect 8582 2942 8612 2957
rect 8683 2942 8713 2957
rect 8773 2942 8803 2957
rect 8892 2942 8922 2957
rect 8082 2925 8118 2942
rect 8172 2925 8208 2942
rect 8053 2909 8119 2925
rect 8053 2875 8069 2909
rect 8103 2875 8119 2909
rect 8053 2859 8119 2875
rect 8161 2909 8227 2925
rect 8161 2875 8177 2909
rect 8211 2875 8227 2909
rect 8161 2859 8227 2875
rect 8059 2813 8089 2859
rect 8167 2813 8197 2859
rect 8269 2828 8305 2942
rect 8386 2901 8422 2942
rect 8487 2925 8523 2942
rect 8356 2885 8422 2901
rect 8356 2851 8372 2885
rect 8406 2851 8422 2885
rect 8464 2909 8530 2925
rect 8464 2875 8480 2909
rect 8514 2875 8530 2909
rect 8579 2901 8615 2942
rect 8464 2859 8530 2875
rect 8572 2885 8638 2901
rect 8356 2835 8422 2851
rect 8269 2813 8299 2828
rect 8387 2813 8417 2835
rect 8473 2813 8503 2859
rect 8572 2851 8588 2885
rect 8622 2851 8638 2885
rect 8572 2835 8638 2851
rect 8602 2813 8632 2835
rect 8680 2828 8716 2942
rect 8770 2925 8806 2942
rect 8889 2925 8925 2942
rect 9056 2940 9092 2957
rect 8758 2909 8824 2925
rect 8758 2875 8774 2909
rect 8808 2875 8824 2909
rect 8758 2859 8824 2875
rect 8872 2909 8938 2925
rect 8872 2875 8888 2909
rect 8922 2875 8938 2909
rect 8872 2862 8938 2875
rect 9056 2924 9190 2940
rect 9056 2890 9072 2924
rect 9106 2890 9140 2924
rect 9174 2890 9190 2924
rect 9307 2920 9343 2963
rect 9840 2959 9870 2974
rect 9943 2959 9973 2974
rect 9837 2932 9873 2959
rect 9056 2874 9190 2890
rect 9238 2904 9343 2920
rect 8680 2813 8710 2828
rect 8766 2813 8796 2859
rect 8872 2832 9008 2862
rect 8978 2813 9008 2832
rect 9123 2813 9153 2874
rect 9238 2870 9254 2904
rect 9288 2870 9343 2904
rect 9238 2854 9343 2870
rect 9825 2916 9891 2932
rect 9940 2916 9976 2959
rect 10041 2949 10077 2980
rect 10449 3153 10479 3179
rect 10550 3153 10580 3179
rect 10642 3153 10672 3179
rect 10740 3168 10776 3221
rect 11116 3183 11152 3221
rect 11370 3198 11400 3224
rect 10743 3153 10773 3168
rect 10833 3153 10863 3179
rect 10952 3153 10982 3179
rect 11119 3168 11149 3183
rect 11902 3194 11932 3220
rect 12103 3217 13214 3247
rect 12103 3206 12139 3217
rect 11119 2953 11149 2968
rect 11370 2959 11400 2974
rect 12005 3170 12035 3196
rect 12106 3191 12136 3206
rect 12207 3149 12237 3175
rect 12297 3149 12327 3175
rect 12391 3164 12427 3217
rect 12394 3149 12424 3164
rect 12106 2976 12136 2991
rect 9825 2882 9841 2916
rect 9875 2882 9891 2916
rect 9825 2866 9891 2882
rect 9933 2900 9999 2916
rect 9933 2866 9949 2900
rect 9983 2866 9999 2900
rect 9313 2832 9343 2854
rect 7780 2658 7810 2684
rect 7903 2659 7933 2685
rect 7981 2659 8011 2685
rect 8059 2659 8089 2685
rect 8167 2659 8197 2685
rect 8269 2659 8299 2685
rect 8387 2659 8417 2685
rect 8473 2659 8503 2685
rect 8602 2659 8632 2685
rect 8680 2659 8710 2685
rect 8766 2659 8796 2685
rect 8978 2659 9008 2685
rect 9123 2659 9153 2685
rect 9840 2828 9870 2866
rect 9933 2850 9999 2866
rect 9313 2658 9343 2684
rect 9963 2809 9993 2850
rect 10041 2809 10071 2949
rect 10145 2938 10175 2953
rect 10235 2938 10265 2953
rect 10332 2938 10362 2953
rect 10449 2938 10479 2953
rect 10550 2938 10580 2953
rect 10642 2938 10672 2953
rect 10743 2938 10773 2953
rect 10833 2938 10863 2953
rect 10952 2938 10982 2953
rect 10142 2921 10178 2938
rect 10232 2921 10268 2938
rect 10113 2905 10179 2921
rect 10113 2871 10129 2905
rect 10163 2871 10179 2905
rect 10113 2855 10179 2871
rect 10221 2905 10287 2921
rect 10221 2871 10237 2905
rect 10271 2871 10287 2905
rect 10221 2855 10287 2871
rect 10119 2809 10149 2855
rect 10227 2809 10257 2855
rect 10329 2824 10365 2938
rect 10446 2897 10482 2938
rect 10547 2921 10583 2938
rect 10416 2881 10482 2897
rect 10416 2847 10432 2881
rect 10466 2847 10482 2881
rect 10524 2905 10590 2921
rect 10524 2871 10540 2905
rect 10574 2871 10590 2905
rect 10639 2897 10675 2938
rect 10524 2855 10590 2871
rect 10632 2881 10698 2897
rect 10416 2831 10482 2847
rect 10329 2809 10359 2824
rect 10447 2809 10477 2831
rect 10533 2809 10563 2855
rect 10632 2847 10648 2881
rect 10682 2847 10698 2881
rect 10632 2831 10698 2847
rect 10662 2809 10692 2831
rect 10740 2824 10776 2938
rect 10830 2921 10866 2938
rect 10949 2921 10985 2938
rect 11116 2936 11152 2953
rect 10818 2905 10884 2921
rect 10818 2871 10834 2905
rect 10868 2871 10884 2905
rect 10818 2855 10884 2871
rect 10932 2905 10998 2921
rect 10932 2871 10948 2905
rect 10982 2871 10998 2905
rect 10932 2858 10998 2871
rect 11116 2920 11250 2936
rect 11116 2886 11132 2920
rect 11166 2886 11200 2920
rect 11234 2886 11250 2920
rect 11367 2916 11403 2959
rect 11902 2955 11932 2970
rect 12005 2955 12035 2970
rect 11899 2928 11935 2955
rect 11116 2870 11250 2886
rect 11298 2900 11403 2916
rect 10740 2809 10770 2824
rect 10826 2809 10856 2855
rect 10932 2828 11068 2858
rect 11038 2809 11068 2828
rect 11183 2809 11213 2870
rect 11298 2866 11314 2900
rect 11348 2866 11403 2900
rect 11298 2850 11403 2866
rect 11887 2912 11953 2928
rect 12002 2912 12038 2955
rect 12103 2945 12139 2976
rect 12511 3149 12541 3175
rect 12612 3149 12642 3175
rect 12704 3149 12734 3175
rect 12802 3164 12838 3217
rect 13178 3179 13214 3217
rect 13432 3194 13462 3220
rect 12805 3149 12835 3164
rect 12895 3149 12925 3175
rect 13014 3149 13044 3175
rect 13181 3164 13211 3179
rect 13976 3192 14006 3218
rect 14177 3215 15288 3245
rect 14177 3204 14213 3215
rect 13181 2949 13211 2964
rect 13432 2955 13462 2970
rect 14079 3168 14109 3194
rect 14180 3189 14210 3204
rect 14281 3147 14311 3173
rect 14371 3147 14401 3173
rect 14465 3162 14501 3215
rect 14468 3147 14498 3162
rect 14180 2974 14210 2989
rect 11887 2878 11903 2912
rect 11937 2878 11953 2912
rect 11887 2862 11953 2878
rect 11995 2896 12061 2912
rect 11995 2862 12011 2896
rect 12045 2862 12061 2896
rect 11373 2828 11403 2850
rect 9840 2654 9870 2680
rect 9963 2655 9993 2681
rect 10041 2655 10071 2681
rect 10119 2655 10149 2681
rect 10227 2655 10257 2681
rect 10329 2655 10359 2681
rect 10447 2655 10477 2681
rect 10533 2655 10563 2681
rect 10662 2655 10692 2681
rect 10740 2655 10770 2681
rect 10826 2655 10856 2681
rect 11038 2655 11068 2681
rect 11183 2655 11213 2681
rect 11902 2824 11932 2862
rect 11995 2846 12061 2862
rect 11373 2654 11403 2680
rect 12025 2805 12055 2846
rect 12103 2805 12133 2945
rect 12207 2934 12237 2949
rect 12297 2934 12327 2949
rect 12394 2934 12424 2949
rect 12511 2934 12541 2949
rect 12612 2934 12642 2949
rect 12704 2934 12734 2949
rect 12805 2934 12835 2949
rect 12895 2934 12925 2949
rect 13014 2934 13044 2949
rect 12204 2917 12240 2934
rect 12294 2917 12330 2934
rect 12175 2901 12241 2917
rect 12175 2867 12191 2901
rect 12225 2867 12241 2901
rect 12175 2851 12241 2867
rect 12283 2901 12349 2917
rect 12283 2867 12299 2901
rect 12333 2867 12349 2901
rect 12283 2851 12349 2867
rect 12181 2805 12211 2851
rect 12289 2805 12319 2851
rect 12391 2820 12427 2934
rect 12508 2893 12544 2934
rect 12609 2917 12645 2934
rect 12478 2877 12544 2893
rect 12478 2843 12494 2877
rect 12528 2843 12544 2877
rect 12586 2901 12652 2917
rect 12586 2867 12602 2901
rect 12636 2867 12652 2901
rect 12701 2893 12737 2934
rect 12586 2851 12652 2867
rect 12694 2877 12760 2893
rect 12478 2827 12544 2843
rect 12391 2805 12421 2820
rect 12509 2805 12539 2827
rect 12595 2805 12625 2851
rect 12694 2843 12710 2877
rect 12744 2843 12760 2877
rect 12694 2827 12760 2843
rect 12724 2805 12754 2827
rect 12802 2820 12838 2934
rect 12892 2917 12928 2934
rect 13011 2917 13047 2934
rect 13178 2932 13214 2949
rect 12880 2901 12946 2917
rect 12880 2867 12896 2901
rect 12930 2867 12946 2901
rect 12880 2851 12946 2867
rect 12994 2901 13060 2917
rect 12994 2867 13010 2901
rect 13044 2867 13060 2901
rect 12994 2854 13060 2867
rect 13178 2916 13312 2932
rect 13178 2882 13194 2916
rect 13228 2882 13262 2916
rect 13296 2882 13312 2916
rect 13429 2912 13465 2955
rect 13976 2953 14006 2968
rect 14079 2953 14109 2968
rect 13973 2926 14009 2953
rect 13178 2866 13312 2882
rect 13360 2896 13465 2912
rect 12802 2805 12832 2820
rect 12888 2805 12918 2851
rect 12994 2824 13130 2854
rect 13100 2805 13130 2824
rect 13245 2805 13275 2866
rect 13360 2862 13376 2896
rect 13410 2862 13465 2896
rect 13360 2846 13465 2862
rect 13961 2910 14027 2926
rect 14076 2910 14112 2953
rect 14177 2943 14213 2974
rect 14585 3147 14615 3173
rect 14686 3147 14716 3173
rect 14778 3147 14808 3173
rect 14876 3162 14912 3215
rect 15252 3177 15288 3215
rect 15506 3192 15536 3218
rect 14879 3147 14909 3162
rect 14969 3147 14999 3173
rect 15088 3147 15118 3173
rect 15255 3162 15285 3177
rect 16038 3188 16068 3214
rect 16239 3211 17350 3241
rect 16239 3200 16275 3211
rect 15255 2947 15285 2962
rect 15506 2953 15536 2968
rect 16141 3164 16171 3190
rect 16242 3185 16272 3200
rect 16343 3143 16373 3169
rect 16433 3143 16463 3169
rect 16527 3158 16563 3211
rect 16530 3143 16560 3158
rect 16242 2970 16272 2985
rect 13961 2876 13977 2910
rect 14011 2876 14027 2910
rect 13961 2860 14027 2876
rect 14069 2894 14135 2910
rect 14069 2860 14085 2894
rect 14119 2860 14135 2894
rect 13435 2824 13465 2846
rect 11902 2650 11932 2676
rect 12025 2651 12055 2677
rect 12103 2651 12133 2677
rect 12181 2651 12211 2677
rect 12289 2651 12319 2677
rect 12391 2651 12421 2677
rect 12509 2651 12539 2677
rect 12595 2651 12625 2677
rect 12724 2651 12754 2677
rect 12802 2651 12832 2677
rect 12888 2651 12918 2677
rect 13100 2651 13130 2677
rect 13245 2651 13275 2677
rect 13976 2822 14006 2860
rect 14069 2844 14135 2860
rect 13435 2650 13465 2676
rect 14099 2803 14129 2844
rect 14177 2803 14207 2943
rect 14281 2932 14311 2947
rect 14371 2932 14401 2947
rect 14468 2932 14498 2947
rect 14585 2932 14615 2947
rect 14686 2932 14716 2947
rect 14778 2932 14808 2947
rect 14879 2932 14909 2947
rect 14969 2932 14999 2947
rect 15088 2932 15118 2947
rect 14278 2915 14314 2932
rect 14368 2915 14404 2932
rect 14249 2899 14315 2915
rect 14249 2865 14265 2899
rect 14299 2865 14315 2899
rect 14249 2849 14315 2865
rect 14357 2899 14423 2915
rect 14357 2865 14373 2899
rect 14407 2865 14423 2899
rect 14357 2849 14423 2865
rect 14255 2803 14285 2849
rect 14363 2803 14393 2849
rect 14465 2818 14501 2932
rect 14582 2891 14618 2932
rect 14683 2915 14719 2932
rect 14552 2875 14618 2891
rect 14552 2841 14568 2875
rect 14602 2841 14618 2875
rect 14660 2899 14726 2915
rect 14660 2865 14676 2899
rect 14710 2865 14726 2899
rect 14775 2891 14811 2932
rect 14660 2849 14726 2865
rect 14768 2875 14834 2891
rect 14552 2825 14618 2841
rect 14465 2803 14495 2818
rect 14583 2803 14613 2825
rect 14669 2803 14699 2849
rect 14768 2841 14784 2875
rect 14818 2841 14834 2875
rect 14768 2825 14834 2841
rect 14798 2803 14828 2825
rect 14876 2818 14912 2932
rect 14966 2915 15002 2932
rect 15085 2915 15121 2932
rect 15252 2930 15288 2947
rect 14954 2899 15020 2915
rect 14954 2865 14970 2899
rect 15004 2865 15020 2899
rect 14954 2849 15020 2865
rect 15068 2899 15134 2915
rect 15068 2865 15084 2899
rect 15118 2865 15134 2899
rect 15068 2852 15134 2865
rect 15252 2914 15386 2930
rect 15252 2880 15268 2914
rect 15302 2880 15336 2914
rect 15370 2880 15386 2914
rect 15503 2910 15539 2953
rect 16038 2949 16068 2964
rect 16141 2949 16171 2964
rect 16035 2922 16071 2949
rect 15252 2864 15386 2880
rect 15434 2894 15539 2910
rect 14876 2803 14906 2818
rect 14962 2803 14992 2849
rect 15068 2822 15204 2852
rect 15174 2803 15204 2822
rect 15319 2803 15349 2864
rect 15434 2860 15450 2894
rect 15484 2860 15539 2894
rect 15434 2844 15539 2860
rect 16023 2906 16089 2922
rect 16138 2906 16174 2949
rect 16239 2939 16275 2970
rect 16647 3143 16677 3169
rect 16748 3143 16778 3169
rect 16840 3143 16870 3169
rect 16938 3158 16974 3211
rect 17314 3173 17350 3211
rect 17568 3188 17598 3214
rect 16941 3143 16971 3158
rect 17031 3143 17061 3169
rect 17150 3143 17180 3169
rect 17317 3158 17347 3173
rect 17317 2943 17347 2958
rect 17568 2949 17598 2964
rect 16023 2872 16039 2906
rect 16073 2872 16089 2906
rect 16023 2856 16089 2872
rect 16131 2890 16197 2906
rect 16131 2856 16147 2890
rect 16181 2856 16197 2890
rect 15509 2822 15539 2844
rect 13976 2648 14006 2674
rect 14099 2649 14129 2675
rect 14177 2649 14207 2675
rect 14255 2649 14285 2675
rect 14363 2649 14393 2675
rect 14465 2649 14495 2675
rect 14583 2649 14613 2675
rect 14669 2649 14699 2675
rect 14798 2649 14828 2675
rect 14876 2649 14906 2675
rect 14962 2649 14992 2675
rect 15174 2649 15204 2675
rect 15319 2649 15349 2675
rect 16038 2818 16068 2856
rect 16131 2840 16197 2856
rect 15509 2648 15539 2674
rect 16161 2799 16191 2840
rect 16239 2799 16269 2939
rect 16343 2928 16373 2943
rect 16433 2928 16463 2943
rect 16530 2928 16560 2943
rect 16647 2928 16677 2943
rect 16748 2928 16778 2943
rect 16840 2928 16870 2943
rect 16941 2928 16971 2943
rect 17031 2928 17061 2943
rect 17150 2928 17180 2943
rect 16340 2911 16376 2928
rect 16430 2911 16466 2928
rect 16311 2895 16377 2911
rect 16311 2861 16327 2895
rect 16361 2861 16377 2895
rect 16311 2845 16377 2861
rect 16419 2895 16485 2911
rect 16419 2861 16435 2895
rect 16469 2861 16485 2895
rect 16419 2845 16485 2861
rect 16317 2799 16347 2845
rect 16425 2799 16455 2845
rect 16527 2814 16563 2928
rect 16644 2887 16680 2928
rect 16745 2911 16781 2928
rect 16614 2871 16680 2887
rect 16614 2837 16630 2871
rect 16664 2837 16680 2871
rect 16722 2895 16788 2911
rect 16722 2861 16738 2895
rect 16772 2861 16788 2895
rect 16837 2887 16873 2928
rect 16722 2845 16788 2861
rect 16830 2871 16896 2887
rect 16614 2821 16680 2837
rect 16527 2799 16557 2814
rect 16645 2799 16675 2821
rect 16731 2799 16761 2845
rect 16830 2837 16846 2871
rect 16880 2837 16896 2871
rect 16830 2821 16896 2837
rect 16860 2799 16890 2821
rect 16938 2814 16974 2928
rect 17028 2911 17064 2928
rect 17147 2911 17183 2928
rect 17314 2926 17350 2943
rect 17016 2895 17082 2911
rect 17016 2861 17032 2895
rect 17066 2861 17082 2895
rect 17016 2845 17082 2861
rect 17130 2895 17196 2911
rect 17130 2861 17146 2895
rect 17180 2861 17196 2895
rect 17130 2848 17196 2861
rect 17314 2910 17448 2926
rect 17314 2876 17330 2910
rect 17364 2876 17398 2910
rect 17432 2876 17448 2910
rect 17565 2906 17601 2949
rect 17314 2860 17448 2876
rect 17496 2890 17601 2906
rect 16938 2799 16968 2814
rect 17024 2799 17054 2845
rect 17130 2818 17266 2848
rect 17236 2799 17266 2818
rect 17381 2799 17411 2860
rect 17496 2856 17512 2890
rect 17546 2856 17601 2890
rect 17496 2840 17601 2856
rect 17571 2818 17601 2840
rect 16038 2644 16068 2670
rect 16161 2645 16191 2671
rect 16239 2645 16269 2671
rect 16317 2645 16347 2671
rect 16425 2645 16455 2671
rect 16527 2645 16557 2671
rect 16645 2645 16675 2671
rect 16731 2645 16761 2671
rect 16860 2645 16890 2671
rect 16938 2645 16968 2671
rect 17024 2645 17054 2671
rect 17236 2645 17266 2671
rect 17381 2645 17411 2671
rect 17571 2644 17601 2670
<< polycont >>
rect 18202 5815 18236 5849
rect 26334 5767 26368 5801
rect 26508 5767 26542 5801
rect 26676 5767 26710 5801
rect 26845 5767 26879 5801
rect 27012 5767 27046 5801
rect 27180 5767 27214 5801
rect 27347 5767 27381 5801
rect 28140 5749 28174 5783
rect 28314 5749 28348 5783
rect 28482 5749 28516 5783
rect 28651 5749 28685 5783
rect 28818 5749 28852 5783
rect 28986 5749 29020 5783
rect 29153 5749 29187 5783
rect 1583 2896 1617 2930
rect 1691 2880 1725 2914
rect 1871 2885 1905 2919
rect 1979 2885 2013 2919
rect 2174 2861 2208 2895
rect 2282 2885 2316 2919
rect 2390 2861 2424 2895
rect 2576 2885 2610 2919
rect 2690 2885 2724 2919
rect 2874 2900 2908 2934
rect 2942 2900 2976 2934
rect 3056 2880 3090 2914
rect 3645 2892 3679 2926
rect 3753 2876 3787 2910
rect 3933 2881 3967 2915
rect 4041 2881 4075 2915
rect 4236 2857 4270 2891
rect 4344 2881 4378 2915
rect 4452 2857 4486 2891
rect 4638 2881 4672 2915
rect 4752 2881 4786 2915
rect 4936 2896 4970 2930
rect 5004 2896 5038 2930
rect 5118 2876 5152 2910
rect 5719 2890 5753 2924
rect 5827 2874 5861 2908
rect 6007 2879 6041 2913
rect 6115 2879 6149 2913
rect 6310 2855 6344 2889
rect 6418 2879 6452 2913
rect 6526 2855 6560 2889
rect 6712 2879 6746 2913
rect 6826 2879 6860 2913
rect 7010 2894 7044 2928
rect 7078 2894 7112 2928
rect 7192 2874 7226 2908
rect 7781 2886 7815 2920
rect 7889 2870 7923 2904
rect 8069 2875 8103 2909
rect 8177 2875 8211 2909
rect 8372 2851 8406 2885
rect 8480 2875 8514 2909
rect 8588 2851 8622 2885
rect 8774 2875 8808 2909
rect 8888 2875 8922 2909
rect 9072 2890 9106 2924
rect 9140 2890 9174 2924
rect 9254 2870 9288 2904
rect 9841 2882 9875 2916
rect 9949 2866 9983 2900
rect 10129 2871 10163 2905
rect 10237 2871 10271 2905
rect 10432 2847 10466 2881
rect 10540 2871 10574 2905
rect 10648 2847 10682 2881
rect 10834 2871 10868 2905
rect 10948 2871 10982 2905
rect 11132 2886 11166 2920
rect 11200 2886 11234 2920
rect 11314 2866 11348 2900
rect 11903 2878 11937 2912
rect 12011 2862 12045 2896
rect 12191 2867 12225 2901
rect 12299 2867 12333 2901
rect 12494 2843 12528 2877
rect 12602 2867 12636 2901
rect 12710 2843 12744 2877
rect 12896 2867 12930 2901
rect 13010 2867 13044 2901
rect 13194 2882 13228 2916
rect 13262 2882 13296 2916
rect 13376 2862 13410 2896
rect 13977 2876 14011 2910
rect 14085 2860 14119 2894
rect 14265 2865 14299 2899
rect 14373 2865 14407 2899
rect 14568 2841 14602 2875
rect 14676 2865 14710 2899
rect 14784 2841 14818 2875
rect 14970 2865 15004 2899
rect 15084 2865 15118 2899
rect 15268 2880 15302 2914
rect 15336 2880 15370 2914
rect 15450 2860 15484 2894
rect 16039 2872 16073 2906
rect 16147 2856 16181 2890
rect 16327 2861 16361 2895
rect 16435 2861 16469 2895
rect 16630 2837 16664 2871
rect 16738 2861 16772 2895
rect 16846 2837 16880 2871
rect 17032 2861 17066 2895
rect 17146 2861 17180 2895
rect 17330 2876 17364 2910
rect 17398 2876 17432 2910
rect 17512 2856 17546 2890
<< locali >>
rect 18122 6127 18151 6161
rect 18185 6127 18243 6161
rect 18277 6127 18335 6161
rect 18369 6127 18398 6161
rect 18190 6085 18232 6127
rect 18190 6051 18198 6085
rect 18190 6017 18232 6051
rect 18190 5983 18198 6017
rect 18190 5949 18232 5983
rect 18190 5915 18198 5949
rect 18190 5899 18232 5915
rect 18266 6085 18332 6093
rect 18266 6051 18282 6085
rect 18316 6051 18332 6085
rect 26292 6079 26321 6113
rect 26355 6079 26413 6113
rect 26447 6079 26505 6113
rect 26539 6079 26597 6113
rect 26631 6079 26689 6113
rect 26723 6079 26781 6113
rect 26815 6079 26873 6113
rect 26907 6079 26965 6113
rect 26999 6079 27057 6113
rect 27091 6079 27149 6113
rect 27183 6079 27241 6113
rect 27275 6079 27333 6113
rect 27367 6079 27425 6113
rect 27459 6079 27517 6113
rect 27551 6079 27609 6113
rect 27643 6079 27701 6113
rect 27735 6079 27764 6113
rect 18266 6017 18332 6051
rect 18266 5983 18282 6017
rect 18316 5983 18332 6017
rect 18266 5949 18332 5983
rect 18266 5915 18282 5949
rect 18316 5915 18332 5949
rect 18266 5897 18332 5915
rect 18186 5854 18252 5863
rect 18186 5816 18196 5854
rect 18186 5815 18202 5816
rect 18236 5815 18252 5854
rect 18286 5852 18332 5897
rect 18286 5818 18298 5852
rect 26332 6037 26374 6079
rect 26332 6003 26340 6037
rect 26332 5969 26374 6003
rect 26332 5935 26340 5969
rect 26332 5899 26374 5935
rect 26332 5865 26340 5899
rect 26332 5849 26374 5865
rect 26408 6037 26474 6045
rect 26408 6003 26424 6037
rect 26458 6003 26474 6037
rect 26408 5969 26474 6003
rect 26408 5935 26424 5969
rect 26458 5935 26474 5969
rect 26408 5899 26474 5935
rect 26508 6037 26542 6079
rect 26508 5969 26542 6003
rect 26508 5919 26542 5935
rect 26576 6037 26642 6045
rect 26576 6003 26592 6037
rect 26626 6003 26642 6037
rect 26576 5969 26642 6003
rect 26576 5935 26592 5969
rect 26626 5935 26642 5969
rect 26408 5865 26424 5899
rect 26458 5885 26474 5899
rect 26576 5899 26642 5935
rect 26676 6037 26710 6079
rect 26676 5969 26710 6003
rect 26676 5919 26710 5935
rect 26744 6037 26810 6045
rect 26744 6003 26760 6037
rect 26794 6003 26810 6037
rect 26744 5969 26810 6003
rect 26744 5935 26760 5969
rect 26794 5935 26810 5969
rect 26576 5885 26592 5899
rect 26458 5865 26592 5885
rect 26626 5885 26642 5899
rect 26744 5899 26810 5935
rect 26844 6037 26878 6079
rect 26844 5969 26878 6003
rect 26844 5919 26878 5935
rect 26912 6037 26978 6045
rect 26912 6003 26928 6037
rect 26962 6003 26978 6037
rect 26912 5969 26978 6003
rect 26912 5935 26928 5969
rect 26962 5935 26978 5969
rect 26744 5885 26760 5899
rect 26626 5865 26760 5885
rect 26794 5885 26810 5899
rect 26912 5899 26978 5935
rect 27012 6037 27046 6079
rect 27012 5969 27046 6003
rect 27012 5919 27046 5935
rect 27080 6037 27146 6045
rect 27080 6003 27096 6037
rect 27130 6003 27146 6037
rect 27080 5969 27146 6003
rect 27080 5935 27096 5969
rect 27130 5935 27146 5969
rect 26912 5885 26928 5899
rect 26794 5865 26928 5885
rect 26962 5885 26978 5899
rect 27080 5899 27146 5935
rect 27180 6037 27214 6079
rect 27180 5969 27214 6003
rect 27180 5919 27214 5935
rect 27248 6037 27314 6045
rect 27248 6003 27264 6037
rect 27298 6003 27314 6037
rect 27248 5969 27314 6003
rect 27248 5935 27264 5969
rect 27298 5935 27314 5969
rect 27080 5885 27096 5899
rect 26962 5865 27096 5885
rect 27130 5885 27146 5899
rect 27248 5899 27314 5935
rect 27348 6037 27382 6079
rect 27348 5969 27382 6003
rect 27348 5919 27382 5935
rect 27416 6037 27482 6045
rect 27416 6003 27432 6037
rect 27466 6003 27482 6037
rect 27416 5969 27482 6003
rect 27416 5935 27432 5969
rect 27466 5935 27482 5969
rect 27248 5885 27264 5899
rect 27130 5865 27264 5885
rect 27298 5885 27314 5899
rect 27416 5899 27482 5935
rect 27516 6037 27550 6079
rect 27516 5969 27550 6003
rect 27516 5919 27550 5935
rect 27584 6037 27650 6045
rect 27584 6003 27600 6037
rect 27634 6003 27650 6037
rect 27584 5969 27650 6003
rect 27584 5935 27600 5969
rect 27634 5935 27650 5969
rect 27416 5885 27432 5899
rect 27298 5865 27432 5885
rect 27466 5885 27482 5899
rect 27584 5899 27650 5935
rect 27684 6037 27726 6079
rect 28098 6061 28127 6095
rect 28161 6061 28219 6095
rect 28253 6061 28311 6095
rect 28345 6061 28403 6095
rect 28437 6061 28495 6095
rect 28529 6061 28587 6095
rect 28621 6061 28679 6095
rect 28713 6061 28771 6095
rect 28805 6061 28863 6095
rect 28897 6061 28955 6095
rect 28989 6061 29047 6095
rect 29081 6061 29139 6095
rect 29173 6061 29231 6095
rect 29265 6061 29323 6095
rect 29357 6061 29415 6095
rect 29449 6061 29507 6095
rect 29541 6061 29570 6095
rect 27718 6003 27726 6037
rect 27684 5969 27726 6003
rect 27718 5935 27726 5969
rect 27684 5919 27726 5935
rect 28138 6019 28180 6061
rect 28138 5985 28146 6019
rect 28138 5951 28180 5985
rect 27584 5885 27600 5899
rect 27466 5865 27600 5885
rect 27634 5865 27650 5899
rect 26408 5851 27650 5865
rect 18186 5765 18232 5781
rect 18286 5777 18332 5818
rect 18186 5731 18198 5765
rect 18186 5697 18232 5731
rect 18186 5663 18198 5697
rect 18186 5617 18232 5663
rect 18266 5765 18332 5777
rect 26309 5810 27397 5815
rect 26309 5801 26364 5810
rect 26406 5801 27397 5810
rect 26309 5767 26334 5801
rect 26406 5772 26508 5801
rect 26368 5767 26508 5772
rect 26542 5767 26676 5801
rect 26710 5767 26845 5801
rect 26879 5767 27012 5801
rect 27046 5767 27180 5801
rect 27214 5767 27347 5801
rect 27381 5767 27397 5801
rect 27584 5794 27650 5851
rect 28138 5917 28146 5951
rect 28138 5881 28180 5917
rect 28138 5847 28146 5881
rect 28138 5831 28180 5847
rect 28214 6019 28280 6027
rect 28214 5985 28230 6019
rect 28264 5985 28280 6019
rect 28214 5951 28280 5985
rect 28214 5917 28230 5951
rect 28264 5917 28280 5951
rect 28214 5881 28280 5917
rect 28314 6019 28348 6061
rect 28314 5951 28348 5985
rect 28314 5901 28348 5917
rect 28382 6019 28448 6027
rect 28382 5985 28398 6019
rect 28432 5985 28448 6019
rect 28382 5951 28448 5985
rect 28382 5917 28398 5951
rect 28432 5917 28448 5951
rect 28214 5847 28230 5881
rect 28264 5867 28280 5881
rect 28382 5881 28448 5917
rect 28482 6019 28516 6061
rect 28482 5951 28516 5985
rect 28482 5901 28516 5917
rect 28550 6019 28616 6027
rect 28550 5985 28566 6019
rect 28600 5985 28616 6019
rect 28550 5951 28616 5985
rect 28550 5917 28566 5951
rect 28600 5917 28616 5951
rect 28382 5867 28398 5881
rect 28264 5847 28398 5867
rect 28432 5867 28448 5881
rect 28550 5881 28616 5917
rect 28650 6019 28684 6061
rect 28650 5951 28684 5985
rect 28650 5901 28684 5917
rect 28718 6019 28784 6027
rect 28718 5985 28734 6019
rect 28768 5985 28784 6019
rect 28718 5951 28784 5985
rect 28718 5917 28734 5951
rect 28768 5917 28784 5951
rect 28550 5867 28566 5881
rect 28432 5847 28566 5867
rect 28600 5867 28616 5881
rect 28718 5881 28784 5917
rect 28818 6019 28852 6061
rect 28818 5951 28852 5985
rect 28818 5901 28852 5917
rect 28886 6019 28952 6027
rect 28886 5985 28902 6019
rect 28936 5985 28952 6019
rect 28886 5951 28952 5985
rect 28886 5917 28902 5951
rect 28936 5917 28952 5951
rect 28718 5867 28734 5881
rect 28600 5847 28734 5867
rect 28768 5867 28784 5881
rect 28886 5881 28952 5917
rect 28986 6019 29020 6061
rect 28986 5951 29020 5985
rect 28986 5901 29020 5917
rect 29054 6019 29120 6027
rect 29054 5985 29070 6019
rect 29104 5985 29120 6019
rect 29054 5951 29120 5985
rect 29054 5917 29070 5951
rect 29104 5917 29120 5951
rect 28886 5867 28902 5881
rect 28768 5847 28902 5867
rect 28936 5867 28952 5881
rect 29054 5881 29120 5917
rect 29154 6019 29188 6061
rect 29154 5951 29188 5985
rect 29154 5901 29188 5917
rect 29222 6019 29288 6027
rect 29222 5985 29238 6019
rect 29272 5985 29288 6019
rect 29222 5951 29288 5985
rect 29222 5917 29238 5951
rect 29272 5917 29288 5951
rect 29054 5867 29070 5881
rect 28936 5847 29070 5867
rect 29104 5867 29120 5881
rect 29222 5881 29288 5917
rect 29322 6019 29356 6061
rect 29322 5951 29356 5985
rect 29322 5901 29356 5917
rect 29390 6019 29456 6027
rect 29390 5985 29406 6019
rect 29440 5985 29456 6019
rect 29390 5951 29456 5985
rect 29390 5917 29406 5951
rect 29440 5917 29456 5951
rect 29222 5867 29238 5881
rect 29104 5847 29238 5867
rect 29272 5867 29288 5881
rect 29390 5881 29456 5917
rect 29490 6019 29532 6061
rect 29524 5985 29532 6019
rect 29490 5951 29532 5985
rect 29524 5917 29532 5951
rect 29490 5901 29532 5917
rect 29390 5867 29406 5881
rect 29272 5847 29406 5867
rect 29440 5847 29456 5881
rect 28214 5833 29456 5847
rect 18266 5731 18282 5765
rect 18316 5731 18332 5765
rect 27584 5756 27600 5794
rect 27640 5756 27650 5794
rect 27584 5733 27650 5756
rect 28115 5792 29203 5797
rect 28115 5783 28170 5792
rect 28212 5783 29203 5792
rect 28115 5749 28140 5783
rect 28212 5754 28314 5783
rect 28174 5749 28314 5754
rect 28348 5749 28482 5783
rect 28516 5749 28651 5783
rect 28685 5749 28818 5783
rect 28852 5749 28986 5783
rect 29020 5749 29153 5783
rect 29187 5749 29203 5783
rect 29390 5776 29456 5833
rect 18266 5697 18332 5731
rect 18266 5663 18282 5697
rect 18316 5663 18332 5697
rect 18266 5651 18332 5663
rect 26328 5713 26374 5729
rect 26328 5679 26340 5713
rect 26328 5645 26374 5679
rect 18122 5583 18151 5617
rect 18185 5583 18243 5617
rect 18277 5583 18335 5617
rect 18369 5583 18398 5617
rect 26328 5611 26340 5645
rect 26328 5569 26374 5611
rect 26408 5713 27650 5733
rect 29390 5738 29406 5776
rect 29446 5738 29456 5776
rect 26408 5679 26424 5713
rect 26458 5695 26592 5713
rect 26458 5679 26474 5695
rect 26408 5645 26474 5679
rect 26576 5679 26592 5695
rect 26626 5695 26760 5713
rect 26626 5679 26642 5695
rect 26408 5611 26424 5645
rect 26458 5611 26474 5645
rect 26408 5603 26474 5611
rect 26508 5645 26542 5661
rect 26508 5569 26542 5611
rect 26576 5645 26642 5679
rect 26744 5679 26760 5695
rect 26794 5695 26928 5713
rect 26794 5679 26810 5695
rect 26576 5611 26592 5645
rect 26626 5611 26642 5645
rect 26576 5603 26642 5611
rect 26676 5645 26710 5661
rect 26676 5569 26710 5611
rect 26744 5645 26810 5679
rect 26912 5679 26928 5695
rect 26962 5695 27096 5713
rect 26962 5679 26978 5695
rect 26744 5611 26760 5645
rect 26794 5611 26810 5645
rect 26744 5603 26810 5611
rect 26844 5645 26878 5661
rect 26844 5569 26878 5611
rect 26912 5645 26978 5679
rect 27080 5679 27096 5695
rect 27130 5695 27264 5713
rect 27130 5679 27146 5695
rect 26912 5611 26928 5645
rect 26962 5611 26978 5645
rect 26912 5603 26978 5611
rect 27012 5645 27046 5661
rect 27012 5569 27046 5611
rect 27080 5645 27146 5679
rect 27248 5679 27264 5695
rect 27298 5695 27432 5713
rect 27298 5679 27314 5695
rect 27080 5611 27096 5645
rect 27130 5611 27146 5645
rect 27080 5603 27146 5611
rect 27180 5645 27214 5661
rect 27180 5569 27214 5611
rect 27248 5645 27314 5679
rect 27416 5679 27432 5695
rect 27466 5695 27600 5713
rect 27466 5679 27482 5695
rect 27248 5611 27264 5645
rect 27298 5611 27314 5645
rect 27248 5603 27314 5611
rect 27348 5645 27382 5661
rect 27348 5569 27382 5611
rect 27416 5645 27482 5679
rect 27584 5679 27600 5695
rect 27634 5679 27650 5713
rect 27416 5611 27432 5645
rect 27466 5611 27482 5645
rect 27416 5603 27482 5611
rect 27516 5645 27550 5661
rect 27516 5569 27550 5611
rect 27584 5645 27650 5679
rect 27584 5611 27600 5645
rect 27634 5611 27650 5645
rect 27584 5603 27650 5611
rect 27684 5713 27726 5729
rect 29390 5715 29456 5738
rect 27718 5679 27726 5713
rect 27684 5645 27726 5679
rect 27718 5611 27726 5645
rect 27684 5569 27726 5611
rect 28134 5695 28180 5711
rect 28134 5661 28146 5695
rect 28134 5627 28180 5661
rect 28134 5593 28146 5627
rect 26292 5535 26321 5569
rect 26355 5535 26413 5569
rect 26447 5535 26505 5569
rect 26539 5535 26597 5569
rect 26631 5535 26689 5569
rect 26723 5535 26781 5569
rect 26815 5535 26873 5569
rect 26907 5535 26965 5569
rect 26999 5535 27057 5569
rect 27091 5535 27149 5569
rect 27183 5535 27241 5569
rect 27275 5535 27333 5569
rect 27367 5535 27425 5569
rect 27459 5535 27517 5569
rect 27551 5535 27609 5569
rect 27643 5535 27701 5569
rect 27735 5535 27764 5569
rect 28134 5551 28180 5593
rect 28214 5695 29456 5715
rect 28214 5661 28230 5695
rect 28264 5677 28398 5695
rect 28264 5661 28280 5677
rect 28214 5627 28280 5661
rect 28382 5661 28398 5677
rect 28432 5677 28566 5695
rect 28432 5661 28448 5677
rect 28214 5593 28230 5627
rect 28264 5593 28280 5627
rect 28214 5585 28280 5593
rect 28314 5627 28348 5643
rect 28314 5551 28348 5593
rect 28382 5627 28448 5661
rect 28550 5661 28566 5677
rect 28600 5677 28734 5695
rect 28600 5661 28616 5677
rect 28382 5593 28398 5627
rect 28432 5593 28448 5627
rect 28382 5585 28448 5593
rect 28482 5627 28516 5643
rect 28482 5551 28516 5593
rect 28550 5627 28616 5661
rect 28718 5661 28734 5677
rect 28768 5677 28902 5695
rect 28768 5661 28784 5677
rect 28550 5593 28566 5627
rect 28600 5593 28616 5627
rect 28550 5585 28616 5593
rect 28650 5627 28684 5643
rect 28650 5551 28684 5593
rect 28718 5627 28784 5661
rect 28886 5661 28902 5677
rect 28936 5677 29070 5695
rect 28936 5661 28952 5677
rect 28718 5593 28734 5627
rect 28768 5593 28784 5627
rect 28718 5585 28784 5593
rect 28818 5627 28852 5643
rect 28818 5551 28852 5593
rect 28886 5627 28952 5661
rect 29054 5661 29070 5677
rect 29104 5677 29238 5695
rect 29104 5661 29120 5677
rect 28886 5593 28902 5627
rect 28936 5593 28952 5627
rect 28886 5585 28952 5593
rect 28986 5627 29020 5643
rect 28986 5551 29020 5593
rect 29054 5627 29120 5661
rect 29222 5661 29238 5677
rect 29272 5677 29406 5695
rect 29272 5661 29288 5677
rect 29054 5593 29070 5627
rect 29104 5593 29120 5627
rect 29054 5585 29120 5593
rect 29154 5627 29188 5643
rect 29154 5551 29188 5593
rect 29222 5627 29288 5661
rect 29390 5661 29406 5677
rect 29440 5661 29456 5695
rect 29222 5593 29238 5627
rect 29272 5593 29288 5627
rect 29222 5585 29288 5593
rect 29322 5627 29356 5643
rect 29322 5551 29356 5593
rect 29390 5627 29456 5661
rect 29390 5593 29406 5627
rect 29440 5593 29456 5627
rect 29390 5585 29456 5593
rect 29490 5695 29532 5711
rect 29524 5661 29532 5695
rect 29490 5627 29532 5661
rect 29524 5593 29532 5627
rect 29490 5551 29532 5593
rect 28098 5517 28127 5551
rect 28161 5517 28219 5551
rect 28253 5517 28311 5551
rect 28345 5517 28403 5551
rect 28437 5517 28495 5551
rect 28529 5517 28587 5551
rect 28621 5517 28679 5551
rect 28713 5517 28771 5551
rect 28805 5517 28863 5551
rect 28897 5517 28955 5551
rect 28989 5517 29047 5551
rect 29081 5517 29139 5551
rect 29173 5517 29231 5551
rect 29265 5517 29323 5551
rect 29357 5517 29415 5551
rect 29449 5517 29507 5551
rect 29541 5517 29570 5551
rect 1498 3269 1529 3303
rect 1563 3269 1625 3303
rect 1659 3269 1721 3303
rect 1755 3269 1817 3303
rect 1851 3269 1913 3303
rect 1947 3269 2009 3303
rect 2043 3269 2105 3303
rect 2139 3269 2201 3303
rect 2235 3269 2297 3303
rect 2331 3269 2393 3303
rect 2427 3269 2489 3303
rect 2523 3269 2585 3303
rect 2619 3269 2681 3303
rect 2715 3269 2777 3303
rect 2811 3269 2873 3303
rect 2907 3269 2969 3303
rect 3003 3269 3065 3303
rect 3099 3269 3161 3303
rect 3195 3269 3226 3303
rect 1515 3200 1569 3216
rect 1515 3166 1535 3200
rect 1515 3117 1569 3166
rect 1515 3083 1535 3117
rect 1515 3034 1569 3083
rect 1515 3000 1535 3034
rect 1609 3200 1675 3269
rect 1609 3166 1625 3200
rect 1659 3166 1675 3200
rect 2114 3196 2180 3269
rect 1609 3132 1675 3166
rect 1609 3098 1625 3132
rect 1659 3098 1675 3132
rect 1609 3064 1675 3098
rect 1609 3030 1625 3064
rect 1659 3030 1675 3064
rect 1914 3155 1980 3171
rect 1914 3121 1930 3155
rect 1964 3121 1980 3155
rect 1914 3087 1980 3121
rect 1914 3053 1930 3087
rect 1964 3053 1980 3087
rect 1914 3044 1980 3053
rect 1515 2984 1569 3000
rect 1709 3019 1980 3044
rect 1709 3010 1930 3019
rect 1709 2996 1743 3010
rect 1515 2846 1549 2984
rect 1605 2962 1743 2996
rect 1914 2985 1930 3010
rect 1964 2985 1980 3019
rect 2020 3155 2070 3171
rect 2054 3121 2070 3155
rect 2114 3162 2130 3196
rect 2164 3162 2180 3196
rect 2114 3146 2180 3162
rect 2020 3112 2070 3121
rect 2218 3128 2284 3171
rect 2218 3112 2234 3128
rect 2020 3094 2234 3112
rect 2268 3094 2284 3128
rect 2020 3078 2284 3094
rect 2319 3131 2385 3269
rect 2319 3097 2335 3131
rect 2369 3097 2385 3131
rect 2319 3081 2385 3097
rect 2512 3155 2597 3171
rect 2512 3121 2528 3155
rect 2562 3121 2597 3155
rect 2020 3063 2070 3078
rect 2054 3029 2070 3063
rect 2512 3044 2597 3121
rect 2020 3013 2070 3029
rect 1811 2970 1857 2976
rect 1605 2946 1639 2962
rect 1583 2930 1639 2946
rect 1617 2896 1639 2930
rect 1811 2936 1817 2970
rect 1851 2936 1857 2970
rect 1914 2969 1980 2985
rect 2104 3010 2528 3044
rect 2562 3010 2597 3044
rect 2631 3155 2688 3171
rect 2631 3121 2647 3155
rect 2681 3121 2688 3155
rect 2631 3071 2688 3121
rect 2722 3157 2863 3269
rect 3049 3200 3115 3269
rect 3560 3265 3591 3299
rect 3625 3265 3687 3299
rect 3721 3265 3783 3299
rect 3817 3265 3879 3299
rect 3913 3265 3975 3299
rect 4009 3265 4071 3299
rect 4105 3265 4167 3299
rect 4201 3265 4263 3299
rect 4297 3265 4359 3299
rect 4393 3265 4455 3299
rect 4489 3265 4551 3299
rect 4585 3265 4647 3299
rect 4681 3265 4743 3299
rect 4777 3265 4839 3299
rect 4873 3265 4935 3299
rect 4969 3265 5031 3299
rect 5065 3265 5127 3299
rect 5161 3265 5223 3299
rect 5257 3265 5288 3299
rect 2722 3123 2738 3157
rect 2772 3123 2813 3157
rect 2847 3123 2863 3157
rect 2722 3120 2863 3123
rect 2898 3170 2962 3186
rect 2898 3136 2912 3170
rect 2946 3136 2962 3170
rect 2898 3071 2962 3136
rect 2631 3037 2647 3071
rect 2681 3060 2962 3071
rect 2681 3037 2912 3060
rect 2896 3026 2912 3037
rect 2946 3026 2962 3060
rect 2896 3010 2962 3026
rect 3049 3166 3065 3200
rect 3099 3166 3115 3200
rect 3049 3117 3115 3166
rect 3049 3083 3065 3117
rect 3099 3083 3115 3117
rect 3049 3034 3115 3083
rect 2104 2979 2138 3010
rect 1811 2935 1857 2936
rect 2014 2945 2138 2979
rect 2563 3003 2597 3010
rect 2266 2970 2337 2976
rect 2014 2935 2048 2945
rect 1583 2880 1639 2896
rect 1515 2830 1571 2846
rect 1515 2796 1537 2830
rect 1515 2740 1571 2796
rect 1515 2706 1537 2740
rect 1605 2770 1639 2880
rect 1675 2914 1741 2928
rect 1675 2880 1691 2914
rect 1725 2880 1741 2914
rect 1675 2864 1741 2880
rect 1811 2919 1921 2935
rect 1811 2885 1871 2919
rect 1905 2885 1921 2919
rect 1811 2872 1921 2885
rect 1963 2919 2048 2935
rect 1963 2885 1979 2919
rect 2013 2885 2048 2919
rect 2266 2936 2297 2970
rect 2331 2936 2337 2970
rect 2266 2919 2337 2936
rect 1963 2872 2048 2885
rect 2158 2895 2224 2911
rect 1707 2838 1741 2864
rect 2158 2861 2174 2895
rect 2208 2861 2224 2895
rect 2266 2885 2282 2919
rect 2316 2885 2337 2919
rect 2483 2970 2529 2976
rect 2483 2936 2489 2970
rect 2523 2936 2529 2970
rect 2563 2969 2808 3003
rect 3049 3000 3065 3034
rect 3099 3000 3115 3034
rect 3049 2984 3115 3000
rect 3155 3200 3206 3216
rect 3189 3166 3206 3200
rect 3155 3117 3206 3166
rect 3189 3083 3206 3117
rect 3155 3034 3206 3083
rect 3189 3000 3206 3034
rect 2483 2935 2529 2936
rect 2483 2919 2626 2935
rect 2266 2872 2337 2885
rect 2374 2896 2440 2911
rect 2374 2895 2396 2896
rect 2158 2838 2224 2861
rect 2374 2861 2390 2895
rect 2430 2862 2440 2896
rect 2483 2885 2576 2919
rect 2610 2885 2626 2919
rect 2483 2875 2626 2885
rect 2660 2919 2740 2935
rect 2660 2885 2690 2919
rect 2724 2885 2740 2919
rect 2660 2884 2740 2885
rect 2424 2861 2440 2862
rect 2374 2841 2440 2861
rect 2660 2841 2694 2884
rect 2774 2850 2808 2969
rect 2858 2940 2992 2976
rect 2858 2934 2920 2940
rect 2960 2934 2992 2940
rect 2858 2900 2874 2934
rect 2908 2900 2920 2934
rect 2976 2900 2992 2934
rect 3155 2960 3206 3000
rect 3577 3196 3631 3212
rect 3577 3162 3597 3196
rect 3577 3113 3631 3162
rect 3577 3079 3597 3113
rect 3577 3030 3631 3079
rect 3577 2996 3597 3030
rect 3671 3196 3737 3265
rect 3671 3162 3687 3196
rect 3721 3162 3737 3196
rect 4176 3192 4242 3265
rect 3671 3128 3737 3162
rect 3671 3094 3687 3128
rect 3721 3094 3737 3128
rect 3671 3060 3737 3094
rect 3671 3026 3687 3060
rect 3721 3026 3737 3060
rect 3976 3151 4042 3167
rect 3976 3117 3992 3151
rect 4026 3117 4042 3151
rect 3976 3083 4042 3117
rect 3976 3049 3992 3083
rect 4026 3049 4042 3083
rect 3976 3040 4042 3049
rect 3577 2980 3631 2996
rect 3771 3015 4042 3040
rect 3771 3006 3992 3015
rect 3771 2992 3805 3006
rect 2858 2898 2920 2900
rect 2960 2898 2992 2900
rect 2858 2884 2992 2898
rect 3040 2914 3106 2930
rect 3040 2880 3056 2914
rect 3090 2880 3106 2914
rect 3040 2850 3106 2880
rect 2374 2838 2694 2841
rect 1707 2807 2694 2838
rect 2728 2816 3106 2850
rect 3155 2926 3174 2960
rect 3155 2846 3206 2926
rect 3140 2830 3206 2846
rect 1707 2804 2440 2807
rect 2728 2773 2762 2816
rect 3140 2796 3156 2830
rect 3190 2796 3206 2830
rect 1605 2747 1952 2770
rect 1605 2736 1902 2747
rect 1515 2690 1571 2706
rect 1886 2713 1902 2736
rect 1936 2713 1952 2747
rect 1623 2668 1641 2702
rect 1675 2668 1694 2702
rect 1886 2691 1952 2713
rect 1994 2754 2280 2770
rect 1994 2720 2018 2754
rect 2052 2736 2230 2754
rect 2052 2720 2076 2736
rect 1994 2704 2076 2720
rect 2214 2720 2230 2736
rect 2264 2720 2280 2754
rect 2214 2704 2280 2720
rect 2314 2746 2409 2762
rect 2314 2712 2344 2746
rect 2378 2712 2409 2746
rect 1623 2637 1694 2668
rect 2112 2668 2128 2702
rect 2162 2668 2178 2702
rect 2112 2637 2178 2668
rect 2314 2637 2409 2712
rect 2507 2757 2762 2773
rect 2507 2723 2523 2757
rect 2557 2739 2762 2757
rect 2796 2766 3016 2782
rect 2796 2748 2966 2766
rect 2557 2723 2573 2739
rect 2507 2707 2573 2723
rect 2796 2705 2830 2748
rect 2950 2732 2966 2748
rect 3000 2732 3016 2766
rect 2950 2716 3016 2732
rect 3054 2758 3104 2774
rect 3054 2724 3070 2758
rect 2609 2671 2625 2705
rect 2659 2671 2719 2705
rect 2753 2671 2830 2705
rect 2864 2698 2914 2714
rect 2898 2664 2914 2698
rect 2864 2637 2914 2664
rect 3054 2637 3104 2724
rect 3140 2740 3206 2796
rect 3140 2706 3156 2740
rect 3190 2706 3206 2740
rect 3140 2690 3206 2706
rect 3577 2842 3611 2980
rect 3667 2958 3805 2992
rect 3976 2981 3992 3006
rect 4026 2981 4042 3015
rect 4082 3151 4132 3167
rect 4116 3117 4132 3151
rect 4176 3158 4192 3192
rect 4226 3158 4242 3192
rect 4176 3142 4242 3158
rect 4082 3108 4132 3117
rect 4280 3124 4346 3167
rect 4280 3108 4296 3124
rect 4082 3090 4296 3108
rect 4330 3090 4346 3124
rect 4082 3074 4346 3090
rect 4381 3127 4447 3265
rect 4381 3093 4397 3127
rect 4431 3093 4447 3127
rect 4381 3077 4447 3093
rect 4574 3151 4659 3167
rect 4574 3117 4590 3151
rect 4624 3117 4659 3151
rect 4082 3059 4132 3074
rect 4116 3025 4132 3059
rect 4574 3040 4659 3117
rect 4082 3009 4132 3025
rect 3873 2966 3919 2972
rect 3667 2942 3701 2958
rect 3645 2926 3701 2942
rect 3679 2892 3701 2926
rect 3873 2932 3879 2966
rect 3913 2932 3919 2966
rect 3976 2965 4042 2981
rect 4166 3006 4590 3040
rect 4624 3006 4659 3040
rect 4693 3151 4750 3167
rect 4693 3117 4709 3151
rect 4743 3117 4750 3151
rect 4693 3067 4750 3117
rect 4784 3153 4925 3265
rect 5111 3196 5177 3265
rect 5634 3263 5665 3297
rect 5699 3263 5761 3297
rect 5795 3263 5857 3297
rect 5891 3263 5953 3297
rect 5987 3263 6049 3297
rect 6083 3263 6145 3297
rect 6179 3263 6241 3297
rect 6275 3263 6337 3297
rect 6371 3263 6433 3297
rect 6467 3263 6529 3297
rect 6563 3263 6625 3297
rect 6659 3263 6721 3297
rect 6755 3263 6817 3297
rect 6851 3263 6913 3297
rect 6947 3263 7009 3297
rect 7043 3263 7105 3297
rect 7139 3263 7201 3297
rect 7235 3263 7297 3297
rect 7331 3263 7362 3297
rect 4784 3119 4800 3153
rect 4834 3119 4875 3153
rect 4909 3119 4925 3153
rect 4784 3116 4925 3119
rect 4960 3166 5024 3182
rect 4960 3132 4974 3166
rect 5008 3132 5024 3166
rect 4960 3067 5024 3132
rect 4693 3033 4709 3067
rect 4743 3056 5024 3067
rect 4743 3033 4974 3056
rect 4958 3022 4974 3033
rect 5008 3022 5024 3056
rect 4958 3006 5024 3022
rect 5111 3162 5127 3196
rect 5161 3162 5177 3196
rect 5111 3113 5177 3162
rect 5111 3079 5127 3113
rect 5161 3079 5177 3113
rect 5111 3030 5177 3079
rect 4166 2975 4200 3006
rect 3873 2931 3919 2932
rect 4076 2941 4200 2975
rect 4625 2999 4659 3006
rect 4328 2966 4399 2972
rect 4076 2931 4110 2941
rect 3645 2876 3701 2892
rect 3577 2826 3633 2842
rect 3577 2792 3599 2826
rect 3577 2736 3633 2792
rect 3577 2702 3599 2736
rect 3667 2766 3701 2876
rect 3737 2910 3803 2924
rect 3737 2876 3753 2910
rect 3787 2876 3803 2910
rect 3737 2860 3803 2876
rect 3873 2915 3983 2931
rect 3873 2881 3933 2915
rect 3967 2881 3983 2915
rect 3873 2868 3983 2881
rect 4025 2915 4110 2931
rect 4025 2881 4041 2915
rect 4075 2881 4110 2915
rect 4328 2932 4359 2966
rect 4393 2932 4399 2966
rect 4328 2915 4399 2932
rect 4025 2868 4110 2881
rect 4220 2891 4286 2907
rect 3769 2834 3803 2860
rect 4220 2857 4236 2891
rect 4270 2857 4286 2891
rect 4328 2881 4344 2915
rect 4378 2881 4399 2915
rect 4545 2966 4591 2972
rect 4545 2932 4551 2966
rect 4585 2932 4591 2966
rect 4625 2965 4870 2999
rect 5111 2996 5127 3030
rect 5161 2996 5177 3030
rect 5111 2980 5177 2996
rect 5217 3196 5268 3212
rect 5251 3162 5268 3196
rect 5217 3113 5268 3162
rect 5251 3079 5268 3113
rect 5217 3030 5268 3079
rect 5251 2996 5268 3030
rect 4545 2931 4591 2932
rect 4545 2915 4688 2931
rect 4328 2868 4399 2881
rect 4436 2892 4502 2907
rect 4436 2891 4458 2892
rect 4220 2834 4286 2857
rect 4436 2857 4452 2891
rect 4492 2858 4502 2892
rect 4545 2881 4638 2915
rect 4672 2881 4688 2915
rect 4545 2871 4688 2881
rect 4722 2915 4802 2931
rect 4722 2881 4752 2915
rect 4786 2881 4802 2915
rect 4722 2880 4802 2881
rect 4486 2857 4502 2858
rect 4436 2837 4502 2857
rect 4722 2837 4756 2880
rect 4836 2846 4870 2965
rect 4920 2936 5054 2972
rect 4920 2930 4982 2936
rect 5022 2930 5054 2936
rect 4920 2896 4936 2930
rect 4970 2896 4982 2930
rect 5038 2896 5054 2930
rect 5217 2962 5268 2996
rect 5217 2928 5232 2962
rect 4920 2894 4982 2896
rect 5022 2894 5054 2896
rect 4920 2880 5054 2894
rect 5102 2910 5168 2926
rect 5102 2876 5118 2910
rect 5152 2876 5168 2910
rect 5102 2846 5168 2876
rect 4436 2834 4756 2837
rect 3769 2803 4756 2834
rect 4790 2812 5168 2846
rect 5217 2842 5268 2928
rect 5202 2826 5268 2842
rect 3769 2800 4502 2803
rect 4790 2769 4824 2812
rect 5202 2792 5218 2826
rect 5252 2792 5268 2826
rect 3667 2743 4014 2766
rect 3667 2732 3964 2743
rect 3577 2686 3633 2702
rect 3948 2709 3964 2732
rect 3998 2709 4014 2743
rect 3685 2664 3703 2698
rect 3737 2664 3756 2698
rect 3948 2687 4014 2709
rect 4056 2750 4342 2766
rect 4056 2716 4080 2750
rect 4114 2732 4292 2750
rect 4114 2716 4138 2732
rect 4056 2700 4138 2716
rect 4276 2716 4292 2732
rect 4326 2716 4342 2750
rect 4276 2700 4342 2716
rect 4376 2742 4471 2758
rect 4376 2708 4406 2742
rect 4440 2708 4471 2742
rect 1498 2603 1529 2637
rect 1563 2603 1625 2637
rect 1659 2603 1721 2637
rect 1755 2603 1817 2637
rect 1851 2603 1913 2637
rect 1947 2603 2009 2637
rect 2043 2603 2105 2637
rect 2139 2603 2201 2637
rect 2235 2603 2297 2637
rect 2331 2603 2393 2637
rect 2427 2603 2489 2637
rect 2523 2603 2585 2637
rect 2619 2603 2681 2637
rect 2715 2603 2777 2637
rect 2811 2603 2873 2637
rect 2907 2603 2969 2637
rect 3003 2603 3065 2637
rect 3099 2603 3161 2637
rect 3195 2603 3226 2637
rect 3685 2633 3756 2664
rect 4174 2664 4190 2698
rect 4224 2664 4240 2698
rect 4174 2633 4240 2664
rect 4376 2633 4471 2708
rect 4569 2753 4824 2769
rect 4569 2719 4585 2753
rect 4619 2735 4824 2753
rect 4858 2762 5078 2778
rect 4858 2744 5028 2762
rect 4619 2719 4635 2735
rect 4569 2703 4635 2719
rect 4858 2701 4892 2744
rect 5012 2728 5028 2744
rect 5062 2728 5078 2762
rect 5012 2712 5078 2728
rect 5116 2754 5166 2770
rect 5116 2720 5132 2754
rect 4671 2667 4687 2701
rect 4721 2667 4781 2701
rect 4815 2667 4892 2701
rect 4926 2694 4976 2710
rect 4960 2660 4976 2694
rect 4926 2633 4976 2660
rect 5116 2633 5166 2720
rect 5202 2736 5268 2792
rect 5202 2702 5218 2736
rect 5252 2702 5268 2736
rect 5202 2686 5268 2702
rect 5651 3194 5705 3210
rect 5651 3160 5671 3194
rect 5651 3111 5705 3160
rect 5651 3077 5671 3111
rect 5651 3028 5705 3077
rect 5651 2994 5671 3028
rect 5745 3194 5811 3263
rect 5745 3160 5761 3194
rect 5795 3160 5811 3194
rect 6250 3190 6316 3263
rect 5745 3126 5811 3160
rect 5745 3092 5761 3126
rect 5795 3092 5811 3126
rect 5745 3058 5811 3092
rect 5745 3024 5761 3058
rect 5795 3024 5811 3058
rect 6050 3149 6116 3165
rect 6050 3115 6066 3149
rect 6100 3115 6116 3149
rect 6050 3081 6116 3115
rect 6050 3047 6066 3081
rect 6100 3047 6116 3081
rect 6050 3038 6116 3047
rect 5651 2978 5705 2994
rect 5845 3013 6116 3038
rect 5845 3004 6066 3013
rect 5845 2990 5879 3004
rect 5651 2840 5685 2978
rect 5741 2956 5879 2990
rect 6050 2979 6066 3004
rect 6100 2979 6116 3013
rect 6156 3149 6206 3165
rect 6190 3115 6206 3149
rect 6250 3156 6266 3190
rect 6300 3156 6316 3190
rect 6250 3140 6316 3156
rect 6156 3106 6206 3115
rect 6354 3122 6420 3165
rect 6354 3106 6370 3122
rect 6156 3088 6370 3106
rect 6404 3088 6420 3122
rect 6156 3072 6420 3088
rect 6455 3125 6521 3263
rect 6455 3091 6471 3125
rect 6505 3091 6521 3125
rect 6455 3075 6521 3091
rect 6648 3149 6733 3165
rect 6648 3115 6664 3149
rect 6698 3115 6733 3149
rect 6156 3057 6206 3072
rect 6190 3023 6206 3057
rect 6648 3038 6733 3115
rect 6156 3007 6206 3023
rect 5947 2964 5993 2970
rect 5741 2940 5775 2956
rect 5719 2924 5775 2940
rect 5753 2890 5775 2924
rect 5947 2930 5953 2964
rect 5987 2930 5993 2964
rect 6050 2963 6116 2979
rect 6240 3004 6664 3038
rect 6698 3004 6733 3038
rect 6767 3149 6824 3165
rect 6767 3115 6783 3149
rect 6817 3115 6824 3149
rect 6767 3065 6824 3115
rect 6858 3151 6999 3263
rect 7185 3194 7251 3263
rect 7696 3259 7727 3293
rect 7761 3259 7823 3293
rect 7857 3259 7919 3293
rect 7953 3259 8015 3293
rect 8049 3259 8111 3293
rect 8145 3259 8207 3293
rect 8241 3259 8303 3293
rect 8337 3259 8399 3293
rect 8433 3259 8495 3293
rect 8529 3259 8591 3293
rect 8625 3259 8687 3293
rect 8721 3259 8783 3293
rect 8817 3259 8879 3293
rect 8913 3259 8975 3293
rect 9009 3259 9071 3293
rect 9105 3259 9167 3293
rect 9201 3259 9263 3293
rect 9297 3259 9359 3293
rect 9393 3259 9424 3293
rect 6858 3117 6874 3151
rect 6908 3117 6949 3151
rect 6983 3117 6999 3151
rect 6858 3114 6999 3117
rect 7034 3164 7098 3180
rect 7034 3130 7048 3164
rect 7082 3130 7098 3164
rect 7034 3065 7098 3130
rect 6767 3031 6783 3065
rect 6817 3054 7098 3065
rect 6817 3031 7048 3054
rect 7032 3020 7048 3031
rect 7082 3020 7098 3054
rect 7032 3004 7098 3020
rect 7185 3160 7201 3194
rect 7235 3160 7251 3194
rect 7185 3111 7251 3160
rect 7185 3077 7201 3111
rect 7235 3077 7251 3111
rect 7185 3028 7251 3077
rect 6240 2973 6274 3004
rect 5947 2929 5993 2930
rect 6150 2939 6274 2973
rect 6699 2997 6733 3004
rect 6402 2964 6473 2970
rect 6150 2929 6184 2939
rect 5719 2874 5775 2890
rect 5651 2824 5707 2840
rect 5651 2790 5673 2824
rect 5651 2734 5707 2790
rect 5651 2700 5673 2734
rect 5741 2764 5775 2874
rect 5811 2908 5877 2922
rect 5811 2874 5827 2908
rect 5861 2874 5877 2908
rect 5811 2858 5877 2874
rect 5947 2913 6057 2929
rect 5947 2879 6007 2913
rect 6041 2879 6057 2913
rect 5947 2866 6057 2879
rect 6099 2913 6184 2929
rect 6099 2879 6115 2913
rect 6149 2879 6184 2913
rect 6402 2930 6433 2964
rect 6467 2930 6473 2964
rect 6402 2913 6473 2930
rect 6099 2866 6184 2879
rect 6294 2889 6360 2905
rect 5843 2832 5877 2858
rect 6294 2855 6310 2889
rect 6344 2855 6360 2889
rect 6402 2879 6418 2913
rect 6452 2879 6473 2913
rect 6619 2964 6665 2970
rect 6619 2930 6625 2964
rect 6659 2930 6665 2964
rect 6699 2963 6944 2997
rect 7185 2994 7201 3028
rect 7235 2994 7251 3028
rect 7185 2978 7251 2994
rect 7291 3194 7342 3210
rect 7325 3160 7342 3194
rect 7291 3111 7342 3160
rect 7325 3077 7342 3111
rect 7291 3028 7342 3077
rect 7325 2994 7342 3028
rect 6619 2929 6665 2930
rect 6619 2913 6762 2929
rect 6402 2866 6473 2879
rect 6510 2890 6576 2905
rect 6510 2889 6532 2890
rect 6294 2832 6360 2855
rect 6510 2855 6526 2889
rect 6566 2856 6576 2890
rect 6619 2879 6712 2913
rect 6746 2879 6762 2913
rect 6619 2869 6762 2879
rect 6796 2913 6876 2929
rect 6796 2879 6826 2913
rect 6860 2879 6876 2913
rect 6796 2878 6876 2879
rect 6560 2855 6576 2856
rect 6510 2835 6576 2855
rect 6796 2835 6830 2878
rect 6910 2844 6944 2963
rect 6994 2934 7128 2970
rect 6994 2928 7056 2934
rect 7096 2928 7128 2934
rect 6994 2894 7010 2928
rect 7044 2894 7056 2928
rect 7112 2894 7128 2928
rect 7291 2954 7342 2994
rect 7713 3190 7767 3206
rect 7713 3156 7733 3190
rect 7713 3107 7767 3156
rect 7713 3073 7733 3107
rect 7713 3024 7767 3073
rect 7713 2990 7733 3024
rect 7807 3190 7873 3259
rect 7807 3156 7823 3190
rect 7857 3156 7873 3190
rect 8312 3186 8378 3259
rect 7807 3122 7873 3156
rect 7807 3088 7823 3122
rect 7857 3088 7873 3122
rect 7807 3054 7873 3088
rect 7807 3020 7823 3054
rect 7857 3020 7873 3054
rect 8112 3145 8178 3161
rect 8112 3111 8128 3145
rect 8162 3111 8178 3145
rect 8112 3077 8178 3111
rect 8112 3043 8128 3077
rect 8162 3043 8178 3077
rect 8112 3034 8178 3043
rect 7713 2974 7767 2990
rect 7907 3009 8178 3034
rect 7907 3000 8128 3009
rect 7907 2986 7941 3000
rect 6994 2892 7056 2894
rect 7096 2892 7128 2894
rect 6994 2878 7128 2892
rect 7176 2908 7242 2924
rect 7176 2874 7192 2908
rect 7226 2874 7242 2908
rect 7176 2844 7242 2874
rect 6510 2832 6830 2835
rect 5843 2801 6830 2832
rect 6864 2810 7242 2844
rect 7291 2920 7310 2954
rect 7291 2840 7342 2920
rect 7276 2824 7342 2840
rect 5843 2798 6576 2801
rect 6864 2767 6898 2810
rect 7276 2790 7292 2824
rect 7326 2790 7342 2824
rect 5741 2741 6088 2764
rect 5741 2730 6038 2741
rect 5651 2684 5707 2700
rect 6022 2707 6038 2730
rect 6072 2707 6088 2741
rect 5759 2662 5777 2696
rect 5811 2662 5830 2696
rect 6022 2685 6088 2707
rect 6130 2748 6416 2764
rect 6130 2714 6154 2748
rect 6188 2730 6366 2748
rect 6188 2714 6212 2730
rect 6130 2698 6212 2714
rect 6350 2714 6366 2730
rect 6400 2714 6416 2748
rect 6350 2698 6416 2714
rect 6450 2740 6545 2756
rect 6450 2706 6480 2740
rect 6514 2706 6545 2740
rect 3560 2599 3591 2633
rect 3625 2599 3687 2633
rect 3721 2599 3783 2633
rect 3817 2599 3879 2633
rect 3913 2599 3975 2633
rect 4009 2599 4071 2633
rect 4105 2599 4167 2633
rect 4201 2599 4263 2633
rect 4297 2599 4359 2633
rect 4393 2599 4455 2633
rect 4489 2599 4551 2633
rect 4585 2599 4647 2633
rect 4681 2599 4743 2633
rect 4777 2599 4839 2633
rect 4873 2599 4935 2633
rect 4969 2599 5031 2633
rect 5065 2599 5127 2633
rect 5161 2599 5223 2633
rect 5257 2599 5288 2633
rect 5759 2631 5830 2662
rect 6248 2662 6264 2696
rect 6298 2662 6314 2696
rect 6248 2631 6314 2662
rect 6450 2631 6545 2706
rect 6643 2751 6898 2767
rect 6643 2717 6659 2751
rect 6693 2733 6898 2751
rect 6932 2760 7152 2776
rect 6932 2742 7102 2760
rect 6693 2717 6709 2733
rect 6643 2701 6709 2717
rect 6932 2699 6966 2742
rect 7086 2726 7102 2742
rect 7136 2726 7152 2760
rect 7086 2710 7152 2726
rect 7190 2752 7240 2768
rect 7190 2718 7206 2752
rect 6745 2665 6761 2699
rect 6795 2665 6855 2699
rect 6889 2665 6966 2699
rect 7000 2692 7050 2708
rect 7034 2658 7050 2692
rect 7000 2631 7050 2658
rect 7190 2631 7240 2718
rect 7276 2734 7342 2790
rect 7276 2700 7292 2734
rect 7326 2700 7342 2734
rect 7276 2684 7342 2700
rect 7713 2836 7747 2974
rect 7803 2952 7941 2986
rect 8112 2975 8128 3000
rect 8162 2975 8178 3009
rect 8218 3145 8268 3161
rect 8252 3111 8268 3145
rect 8312 3152 8328 3186
rect 8362 3152 8378 3186
rect 8312 3136 8378 3152
rect 8218 3102 8268 3111
rect 8416 3118 8482 3161
rect 8416 3102 8432 3118
rect 8218 3084 8432 3102
rect 8466 3084 8482 3118
rect 8218 3068 8482 3084
rect 8517 3121 8583 3259
rect 8517 3087 8533 3121
rect 8567 3087 8583 3121
rect 8517 3071 8583 3087
rect 8710 3145 8795 3161
rect 8710 3111 8726 3145
rect 8760 3111 8795 3145
rect 8218 3053 8268 3068
rect 8252 3019 8268 3053
rect 8710 3034 8795 3111
rect 8218 3003 8268 3019
rect 8009 2960 8055 2966
rect 7803 2936 7837 2952
rect 7781 2920 7837 2936
rect 7815 2886 7837 2920
rect 8009 2926 8015 2960
rect 8049 2926 8055 2960
rect 8112 2959 8178 2975
rect 8302 3000 8726 3034
rect 8760 3000 8795 3034
rect 8829 3145 8886 3161
rect 8829 3111 8845 3145
rect 8879 3111 8886 3145
rect 8829 3061 8886 3111
rect 8920 3147 9061 3259
rect 9247 3190 9313 3259
rect 9756 3255 9787 3289
rect 9821 3255 9883 3289
rect 9917 3255 9979 3289
rect 10013 3255 10075 3289
rect 10109 3255 10171 3289
rect 10205 3255 10267 3289
rect 10301 3255 10363 3289
rect 10397 3255 10459 3289
rect 10493 3255 10555 3289
rect 10589 3255 10651 3289
rect 10685 3255 10747 3289
rect 10781 3255 10843 3289
rect 10877 3255 10939 3289
rect 10973 3255 11035 3289
rect 11069 3255 11131 3289
rect 11165 3255 11227 3289
rect 11261 3255 11323 3289
rect 11357 3255 11419 3289
rect 11453 3255 11484 3289
rect 8920 3113 8936 3147
rect 8970 3113 9011 3147
rect 9045 3113 9061 3147
rect 8920 3110 9061 3113
rect 9096 3160 9160 3176
rect 9096 3126 9110 3160
rect 9144 3126 9160 3160
rect 9096 3061 9160 3126
rect 8829 3027 8845 3061
rect 8879 3050 9160 3061
rect 8879 3027 9110 3050
rect 9094 3016 9110 3027
rect 9144 3016 9160 3050
rect 9094 3000 9160 3016
rect 9247 3156 9263 3190
rect 9297 3156 9313 3190
rect 9247 3107 9313 3156
rect 9247 3073 9263 3107
rect 9297 3073 9313 3107
rect 9247 3024 9313 3073
rect 8302 2969 8336 3000
rect 8009 2925 8055 2926
rect 8212 2935 8336 2969
rect 8761 2993 8795 3000
rect 8464 2960 8535 2966
rect 8212 2925 8246 2935
rect 7781 2870 7837 2886
rect 7713 2820 7769 2836
rect 7713 2786 7735 2820
rect 7713 2730 7769 2786
rect 7713 2696 7735 2730
rect 7803 2760 7837 2870
rect 7873 2904 7939 2918
rect 7873 2870 7889 2904
rect 7923 2870 7939 2904
rect 7873 2854 7939 2870
rect 8009 2909 8119 2925
rect 8009 2875 8069 2909
rect 8103 2875 8119 2909
rect 8009 2862 8119 2875
rect 8161 2909 8246 2925
rect 8161 2875 8177 2909
rect 8211 2875 8246 2909
rect 8464 2926 8495 2960
rect 8529 2926 8535 2960
rect 8464 2909 8535 2926
rect 8161 2862 8246 2875
rect 8356 2885 8422 2901
rect 7905 2828 7939 2854
rect 8356 2851 8372 2885
rect 8406 2851 8422 2885
rect 8464 2875 8480 2909
rect 8514 2875 8535 2909
rect 8681 2960 8727 2966
rect 8681 2926 8687 2960
rect 8721 2926 8727 2960
rect 8761 2959 9006 2993
rect 9247 2990 9263 3024
rect 9297 2990 9313 3024
rect 9247 2974 9313 2990
rect 9353 3190 9404 3206
rect 9387 3156 9404 3190
rect 9353 3107 9404 3156
rect 9387 3073 9404 3107
rect 9353 3024 9404 3073
rect 9387 2990 9404 3024
rect 8681 2925 8727 2926
rect 8681 2909 8824 2925
rect 8464 2862 8535 2875
rect 8572 2886 8638 2901
rect 8572 2885 8594 2886
rect 8356 2828 8422 2851
rect 8572 2851 8588 2885
rect 8628 2852 8638 2886
rect 8681 2875 8774 2909
rect 8808 2875 8824 2909
rect 8681 2865 8824 2875
rect 8858 2909 8938 2925
rect 8858 2875 8888 2909
rect 8922 2875 8938 2909
rect 8858 2874 8938 2875
rect 8622 2851 8638 2852
rect 8572 2831 8638 2851
rect 8858 2831 8892 2874
rect 8972 2840 9006 2959
rect 9056 2930 9190 2966
rect 9056 2924 9118 2930
rect 9158 2924 9190 2930
rect 9056 2890 9072 2924
rect 9106 2890 9118 2924
rect 9174 2890 9190 2924
rect 9353 2944 9404 2990
rect 9056 2888 9118 2890
rect 9158 2888 9190 2890
rect 9056 2874 9190 2888
rect 9238 2904 9304 2920
rect 9238 2870 9254 2904
rect 9288 2870 9304 2904
rect 9238 2840 9304 2870
rect 8572 2828 8892 2831
rect 7905 2797 8892 2828
rect 8926 2806 9304 2840
rect 9353 2910 9366 2944
rect 9402 2910 9404 2944
rect 9353 2836 9404 2910
rect 9338 2820 9404 2836
rect 7905 2794 8638 2797
rect 8926 2763 8960 2806
rect 9338 2786 9354 2820
rect 9388 2786 9404 2820
rect 7803 2737 8150 2760
rect 7803 2726 8100 2737
rect 7713 2680 7769 2696
rect 8084 2703 8100 2726
rect 8134 2703 8150 2737
rect 7821 2658 7839 2692
rect 7873 2658 7892 2692
rect 8084 2681 8150 2703
rect 8192 2744 8478 2760
rect 8192 2710 8216 2744
rect 8250 2726 8428 2744
rect 8250 2710 8274 2726
rect 8192 2694 8274 2710
rect 8412 2710 8428 2726
rect 8462 2710 8478 2744
rect 8412 2694 8478 2710
rect 8512 2736 8607 2752
rect 8512 2702 8542 2736
rect 8576 2702 8607 2736
rect 5634 2597 5665 2631
rect 5699 2597 5761 2631
rect 5795 2597 5857 2631
rect 5891 2597 5953 2631
rect 5987 2597 6049 2631
rect 6083 2597 6145 2631
rect 6179 2597 6241 2631
rect 6275 2597 6337 2631
rect 6371 2597 6433 2631
rect 6467 2597 6529 2631
rect 6563 2597 6625 2631
rect 6659 2597 6721 2631
rect 6755 2597 6817 2631
rect 6851 2597 6913 2631
rect 6947 2597 7009 2631
rect 7043 2597 7105 2631
rect 7139 2597 7201 2631
rect 7235 2597 7297 2631
rect 7331 2597 7362 2631
rect 7821 2627 7892 2658
rect 8310 2658 8326 2692
rect 8360 2658 8376 2692
rect 8310 2627 8376 2658
rect 8512 2627 8607 2702
rect 8705 2747 8960 2763
rect 8705 2713 8721 2747
rect 8755 2729 8960 2747
rect 8994 2756 9214 2772
rect 8994 2738 9164 2756
rect 8755 2713 8771 2729
rect 8705 2697 8771 2713
rect 8994 2695 9028 2738
rect 9148 2722 9164 2738
rect 9198 2722 9214 2756
rect 9148 2706 9214 2722
rect 9252 2748 9302 2764
rect 9252 2714 9268 2748
rect 8807 2661 8823 2695
rect 8857 2661 8917 2695
rect 8951 2661 9028 2695
rect 9062 2688 9112 2704
rect 9096 2654 9112 2688
rect 9062 2627 9112 2654
rect 9252 2627 9302 2714
rect 9338 2730 9404 2786
rect 9338 2696 9354 2730
rect 9388 2696 9404 2730
rect 9338 2680 9404 2696
rect 9773 3186 9827 3202
rect 9773 3152 9793 3186
rect 9773 3103 9827 3152
rect 9773 3069 9793 3103
rect 9773 3020 9827 3069
rect 9773 2986 9793 3020
rect 9867 3186 9933 3255
rect 9867 3152 9883 3186
rect 9917 3152 9933 3186
rect 10372 3182 10438 3255
rect 9867 3118 9933 3152
rect 9867 3084 9883 3118
rect 9917 3084 9933 3118
rect 9867 3050 9933 3084
rect 9867 3016 9883 3050
rect 9917 3016 9933 3050
rect 10172 3141 10238 3157
rect 10172 3107 10188 3141
rect 10222 3107 10238 3141
rect 10172 3073 10238 3107
rect 10172 3039 10188 3073
rect 10222 3039 10238 3073
rect 10172 3030 10238 3039
rect 9773 2970 9827 2986
rect 9967 3005 10238 3030
rect 9967 2996 10188 3005
rect 9967 2982 10001 2996
rect 9773 2832 9807 2970
rect 9863 2948 10001 2982
rect 10172 2971 10188 2996
rect 10222 2971 10238 3005
rect 10278 3141 10328 3157
rect 10312 3107 10328 3141
rect 10372 3148 10388 3182
rect 10422 3148 10438 3182
rect 10372 3132 10438 3148
rect 10278 3098 10328 3107
rect 10476 3114 10542 3157
rect 10476 3098 10492 3114
rect 10278 3080 10492 3098
rect 10526 3080 10542 3114
rect 10278 3064 10542 3080
rect 10577 3117 10643 3255
rect 10577 3083 10593 3117
rect 10627 3083 10643 3117
rect 10577 3067 10643 3083
rect 10770 3141 10855 3157
rect 10770 3107 10786 3141
rect 10820 3107 10855 3141
rect 10278 3049 10328 3064
rect 10312 3015 10328 3049
rect 10770 3030 10855 3107
rect 10278 2999 10328 3015
rect 10069 2956 10115 2962
rect 9863 2932 9897 2948
rect 9841 2916 9897 2932
rect 9875 2882 9897 2916
rect 10069 2922 10075 2956
rect 10109 2922 10115 2956
rect 10172 2955 10238 2971
rect 10362 2996 10786 3030
rect 10820 2996 10855 3030
rect 10889 3141 10946 3157
rect 10889 3107 10905 3141
rect 10939 3107 10946 3141
rect 10889 3057 10946 3107
rect 10980 3143 11121 3255
rect 11307 3186 11373 3255
rect 11818 3251 11849 3285
rect 11883 3251 11945 3285
rect 11979 3251 12041 3285
rect 12075 3251 12137 3285
rect 12171 3251 12233 3285
rect 12267 3251 12329 3285
rect 12363 3251 12425 3285
rect 12459 3251 12521 3285
rect 12555 3251 12617 3285
rect 12651 3251 12713 3285
rect 12747 3251 12809 3285
rect 12843 3251 12905 3285
rect 12939 3251 13001 3285
rect 13035 3251 13097 3285
rect 13131 3251 13193 3285
rect 13227 3251 13289 3285
rect 13323 3251 13385 3285
rect 13419 3251 13481 3285
rect 13515 3251 13546 3285
rect 10980 3109 10996 3143
rect 11030 3109 11071 3143
rect 11105 3109 11121 3143
rect 10980 3106 11121 3109
rect 11156 3156 11220 3172
rect 11156 3122 11170 3156
rect 11204 3122 11220 3156
rect 11156 3057 11220 3122
rect 10889 3023 10905 3057
rect 10939 3046 11220 3057
rect 10939 3023 11170 3046
rect 11154 3012 11170 3023
rect 11204 3012 11220 3046
rect 11154 2996 11220 3012
rect 11307 3152 11323 3186
rect 11357 3152 11373 3186
rect 11307 3103 11373 3152
rect 11307 3069 11323 3103
rect 11357 3069 11373 3103
rect 11307 3020 11373 3069
rect 10362 2965 10396 2996
rect 10069 2921 10115 2922
rect 10272 2931 10396 2965
rect 10821 2989 10855 2996
rect 10524 2956 10595 2962
rect 10272 2921 10306 2931
rect 9841 2866 9897 2882
rect 9773 2816 9829 2832
rect 9773 2782 9795 2816
rect 9773 2726 9829 2782
rect 9773 2692 9795 2726
rect 9863 2756 9897 2866
rect 9933 2900 9999 2914
rect 9933 2866 9949 2900
rect 9983 2866 9999 2900
rect 9933 2850 9999 2866
rect 10069 2905 10179 2921
rect 10069 2871 10129 2905
rect 10163 2871 10179 2905
rect 10069 2858 10179 2871
rect 10221 2905 10306 2921
rect 10221 2871 10237 2905
rect 10271 2871 10306 2905
rect 10524 2922 10555 2956
rect 10589 2922 10595 2956
rect 10524 2905 10595 2922
rect 10221 2858 10306 2871
rect 10416 2881 10482 2897
rect 9965 2824 9999 2850
rect 10416 2847 10432 2881
rect 10466 2847 10482 2881
rect 10524 2871 10540 2905
rect 10574 2871 10595 2905
rect 10741 2956 10787 2962
rect 10741 2922 10747 2956
rect 10781 2922 10787 2956
rect 10821 2955 11066 2989
rect 11307 2986 11323 3020
rect 11357 2986 11373 3020
rect 11307 2970 11373 2986
rect 11413 3186 11464 3202
rect 11447 3152 11464 3186
rect 11413 3103 11464 3152
rect 11447 3069 11464 3103
rect 11413 3020 11464 3069
rect 11447 2986 11464 3020
rect 10741 2921 10787 2922
rect 10741 2905 10884 2921
rect 10524 2858 10595 2871
rect 10632 2882 10698 2897
rect 10632 2881 10654 2882
rect 10416 2824 10482 2847
rect 10632 2847 10648 2881
rect 10688 2848 10698 2882
rect 10741 2871 10834 2905
rect 10868 2871 10884 2905
rect 10741 2861 10884 2871
rect 10918 2905 10998 2921
rect 10918 2871 10948 2905
rect 10982 2871 10998 2905
rect 10918 2870 10998 2871
rect 10682 2847 10698 2848
rect 10632 2827 10698 2847
rect 10918 2827 10952 2870
rect 11032 2836 11066 2955
rect 11116 2926 11250 2962
rect 11116 2920 11178 2926
rect 11218 2920 11250 2926
rect 11116 2886 11132 2920
rect 11166 2886 11178 2920
rect 11234 2886 11250 2920
rect 11413 2946 11464 2986
rect 11835 3182 11889 3198
rect 11835 3148 11855 3182
rect 11835 3099 11889 3148
rect 11835 3065 11855 3099
rect 11835 3016 11889 3065
rect 11835 2982 11855 3016
rect 11929 3182 11995 3251
rect 11929 3148 11945 3182
rect 11979 3148 11995 3182
rect 12434 3178 12500 3251
rect 11929 3114 11995 3148
rect 11929 3080 11945 3114
rect 11979 3080 11995 3114
rect 11929 3046 11995 3080
rect 11929 3012 11945 3046
rect 11979 3012 11995 3046
rect 12234 3137 12300 3153
rect 12234 3103 12250 3137
rect 12284 3103 12300 3137
rect 12234 3069 12300 3103
rect 12234 3035 12250 3069
rect 12284 3035 12300 3069
rect 12234 3026 12300 3035
rect 11835 2966 11889 2982
rect 12029 3001 12300 3026
rect 12029 2992 12250 3001
rect 12029 2978 12063 2992
rect 11116 2884 11178 2886
rect 11218 2884 11250 2886
rect 11116 2870 11250 2884
rect 11298 2900 11364 2916
rect 11298 2866 11314 2900
rect 11348 2866 11364 2900
rect 11298 2836 11364 2866
rect 10632 2824 10952 2827
rect 9965 2793 10952 2824
rect 10986 2802 11364 2836
rect 11413 2912 11432 2946
rect 11413 2832 11464 2912
rect 11398 2816 11464 2832
rect 9965 2790 10698 2793
rect 10986 2759 11020 2802
rect 11398 2782 11414 2816
rect 11448 2782 11464 2816
rect 9863 2733 10210 2756
rect 9863 2722 10160 2733
rect 9773 2676 9829 2692
rect 10144 2699 10160 2722
rect 10194 2699 10210 2733
rect 9881 2654 9899 2688
rect 9933 2654 9952 2688
rect 10144 2677 10210 2699
rect 10252 2740 10538 2756
rect 10252 2706 10276 2740
rect 10310 2722 10488 2740
rect 10310 2706 10334 2722
rect 10252 2690 10334 2706
rect 10472 2706 10488 2722
rect 10522 2706 10538 2740
rect 10472 2690 10538 2706
rect 10572 2732 10667 2748
rect 10572 2698 10602 2732
rect 10636 2698 10667 2732
rect 7696 2593 7727 2627
rect 7761 2593 7823 2627
rect 7857 2593 7919 2627
rect 7953 2593 8015 2627
rect 8049 2593 8111 2627
rect 8145 2593 8207 2627
rect 8241 2593 8303 2627
rect 8337 2593 8399 2627
rect 8433 2593 8495 2627
rect 8529 2593 8591 2627
rect 8625 2593 8687 2627
rect 8721 2593 8783 2627
rect 8817 2593 8879 2627
rect 8913 2593 8975 2627
rect 9009 2593 9071 2627
rect 9105 2593 9167 2627
rect 9201 2593 9263 2627
rect 9297 2593 9359 2627
rect 9393 2593 9424 2627
rect 9881 2623 9952 2654
rect 10370 2654 10386 2688
rect 10420 2654 10436 2688
rect 10370 2623 10436 2654
rect 10572 2623 10667 2698
rect 10765 2743 11020 2759
rect 10765 2709 10781 2743
rect 10815 2725 11020 2743
rect 11054 2752 11274 2768
rect 11054 2734 11224 2752
rect 10815 2709 10831 2725
rect 10765 2693 10831 2709
rect 11054 2691 11088 2734
rect 11208 2718 11224 2734
rect 11258 2718 11274 2752
rect 11208 2702 11274 2718
rect 11312 2744 11362 2760
rect 11312 2710 11328 2744
rect 10867 2657 10883 2691
rect 10917 2657 10977 2691
rect 11011 2657 11088 2691
rect 11122 2684 11172 2700
rect 11156 2650 11172 2684
rect 11122 2623 11172 2650
rect 11312 2623 11362 2710
rect 11398 2726 11464 2782
rect 11398 2692 11414 2726
rect 11448 2692 11464 2726
rect 11398 2676 11464 2692
rect 11835 2828 11869 2966
rect 11925 2944 12063 2978
rect 12234 2967 12250 2992
rect 12284 2967 12300 3001
rect 12340 3137 12390 3153
rect 12374 3103 12390 3137
rect 12434 3144 12450 3178
rect 12484 3144 12500 3178
rect 12434 3128 12500 3144
rect 12340 3094 12390 3103
rect 12538 3110 12604 3153
rect 12538 3094 12554 3110
rect 12340 3076 12554 3094
rect 12588 3076 12604 3110
rect 12340 3060 12604 3076
rect 12639 3113 12705 3251
rect 12639 3079 12655 3113
rect 12689 3079 12705 3113
rect 12639 3063 12705 3079
rect 12832 3137 12917 3153
rect 12832 3103 12848 3137
rect 12882 3103 12917 3137
rect 12340 3045 12390 3060
rect 12374 3011 12390 3045
rect 12832 3026 12917 3103
rect 12340 2995 12390 3011
rect 12131 2952 12177 2958
rect 11925 2928 11959 2944
rect 11903 2912 11959 2928
rect 11937 2878 11959 2912
rect 12131 2918 12137 2952
rect 12171 2918 12177 2952
rect 12234 2951 12300 2967
rect 12424 2992 12848 3026
rect 12882 2992 12917 3026
rect 12951 3137 13008 3153
rect 12951 3103 12967 3137
rect 13001 3103 13008 3137
rect 12951 3053 13008 3103
rect 13042 3139 13183 3251
rect 13369 3182 13435 3251
rect 13892 3249 13923 3283
rect 13957 3249 14019 3283
rect 14053 3249 14115 3283
rect 14149 3249 14211 3283
rect 14245 3249 14307 3283
rect 14341 3249 14403 3283
rect 14437 3249 14499 3283
rect 14533 3249 14595 3283
rect 14629 3249 14691 3283
rect 14725 3249 14787 3283
rect 14821 3249 14883 3283
rect 14917 3249 14979 3283
rect 15013 3249 15075 3283
rect 15109 3249 15171 3283
rect 15205 3249 15267 3283
rect 15301 3249 15363 3283
rect 15397 3249 15459 3283
rect 15493 3249 15555 3283
rect 15589 3249 15620 3283
rect 13042 3105 13058 3139
rect 13092 3105 13133 3139
rect 13167 3105 13183 3139
rect 13042 3102 13183 3105
rect 13218 3152 13282 3168
rect 13218 3118 13232 3152
rect 13266 3118 13282 3152
rect 13218 3053 13282 3118
rect 12951 3019 12967 3053
rect 13001 3042 13282 3053
rect 13001 3019 13232 3042
rect 13216 3008 13232 3019
rect 13266 3008 13282 3042
rect 13216 2992 13282 3008
rect 13369 3148 13385 3182
rect 13419 3148 13435 3182
rect 13369 3099 13435 3148
rect 13369 3065 13385 3099
rect 13419 3065 13435 3099
rect 13369 3016 13435 3065
rect 12424 2961 12458 2992
rect 12131 2917 12177 2918
rect 12334 2927 12458 2961
rect 12883 2985 12917 2992
rect 12586 2952 12657 2958
rect 12334 2917 12368 2927
rect 11903 2862 11959 2878
rect 11835 2812 11891 2828
rect 11835 2778 11857 2812
rect 11835 2722 11891 2778
rect 11835 2688 11857 2722
rect 11925 2752 11959 2862
rect 11995 2896 12061 2910
rect 11995 2862 12011 2896
rect 12045 2862 12061 2896
rect 11995 2846 12061 2862
rect 12131 2901 12241 2917
rect 12131 2867 12191 2901
rect 12225 2867 12241 2901
rect 12131 2854 12241 2867
rect 12283 2901 12368 2917
rect 12283 2867 12299 2901
rect 12333 2867 12368 2901
rect 12586 2918 12617 2952
rect 12651 2918 12657 2952
rect 12586 2901 12657 2918
rect 12283 2854 12368 2867
rect 12478 2877 12544 2893
rect 12027 2820 12061 2846
rect 12478 2843 12494 2877
rect 12528 2843 12544 2877
rect 12586 2867 12602 2901
rect 12636 2867 12657 2901
rect 12803 2952 12849 2958
rect 12803 2918 12809 2952
rect 12843 2918 12849 2952
rect 12883 2951 13128 2985
rect 13369 2982 13385 3016
rect 13419 2982 13435 3016
rect 13369 2966 13435 2982
rect 13475 3182 13526 3198
rect 13509 3148 13526 3182
rect 13475 3099 13526 3148
rect 13509 3065 13526 3099
rect 13475 3016 13526 3065
rect 13509 2982 13526 3016
rect 12803 2917 12849 2918
rect 12803 2901 12946 2917
rect 12586 2854 12657 2867
rect 12694 2878 12760 2893
rect 12694 2877 12716 2878
rect 12478 2820 12544 2843
rect 12694 2843 12710 2877
rect 12750 2844 12760 2878
rect 12803 2867 12896 2901
rect 12930 2867 12946 2901
rect 12803 2857 12946 2867
rect 12980 2901 13060 2917
rect 12980 2867 13010 2901
rect 13044 2867 13060 2901
rect 12980 2866 13060 2867
rect 12744 2843 12760 2844
rect 12694 2823 12760 2843
rect 12980 2823 13014 2866
rect 13094 2832 13128 2951
rect 13178 2922 13312 2958
rect 13178 2916 13240 2922
rect 13280 2916 13312 2922
rect 13178 2882 13194 2916
rect 13228 2882 13240 2916
rect 13296 2882 13312 2916
rect 13475 2948 13526 2982
rect 13475 2914 13490 2948
rect 13178 2880 13240 2882
rect 13280 2880 13312 2882
rect 13178 2866 13312 2880
rect 13360 2896 13426 2912
rect 13360 2862 13376 2896
rect 13410 2862 13426 2896
rect 13360 2832 13426 2862
rect 12694 2820 13014 2823
rect 12027 2789 13014 2820
rect 13048 2798 13426 2832
rect 13475 2828 13526 2914
rect 13460 2812 13526 2828
rect 12027 2786 12760 2789
rect 13048 2755 13082 2798
rect 13460 2778 13476 2812
rect 13510 2778 13526 2812
rect 11925 2729 12272 2752
rect 11925 2718 12222 2729
rect 11835 2672 11891 2688
rect 12206 2695 12222 2718
rect 12256 2695 12272 2729
rect 11943 2650 11961 2684
rect 11995 2650 12014 2684
rect 12206 2673 12272 2695
rect 12314 2736 12600 2752
rect 12314 2702 12338 2736
rect 12372 2718 12550 2736
rect 12372 2702 12396 2718
rect 12314 2686 12396 2702
rect 12534 2702 12550 2718
rect 12584 2702 12600 2736
rect 12534 2686 12600 2702
rect 12634 2728 12729 2744
rect 12634 2694 12664 2728
rect 12698 2694 12729 2728
rect 9756 2589 9787 2623
rect 9821 2589 9883 2623
rect 9917 2589 9979 2623
rect 10013 2589 10075 2623
rect 10109 2589 10171 2623
rect 10205 2589 10267 2623
rect 10301 2589 10363 2623
rect 10397 2589 10459 2623
rect 10493 2589 10555 2623
rect 10589 2589 10651 2623
rect 10685 2589 10747 2623
rect 10781 2589 10843 2623
rect 10877 2589 10939 2623
rect 10973 2589 11035 2623
rect 11069 2589 11131 2623
rect 11165 2589 11227 2623
rect 11261 2589 11323 2623
rect 11357 2589 11419 2623
rect 11453 2589 11484 2623
rect 11943 2619 12014 2650
rect 12432 2650 12448 2684
rect 12482 2650 12498 2684
rect 12432 2619 12498 2650
rect 12634 2619 12729 2694
rect 12827 2739 13082 2755
rect 12827 2705 12843 2739
rect 12877 2721 13082 2739
rect 13116 2748 13336 2764
rect 13116 2730 13286 2748
rect 12877 2705 12893 2721
rect 12827 2689 12893 2705
rect 13116 2687 13150 2730
rect 13270 2714 13286 2730
rect 13320 2714 13336 2748
rect 13270 2698 13336 2714
rect 13374 2740 13424 2756
rect 13374 2706 13390 2740
rect 12929 2653 12945 2687
rect 12979 2653 13039 2687
rect 13073 2653 13150 2687
rect 13184 2680 13234 2696
rect 13218 2646 13234 2680
rect 13184 2619 13234 2646
rect 13374 2619 13424 2706
rect 13460 2722 13526 2778
rect 13460 2688 13476 2722
rect 13510 2688 13526 2722
rect 13460 2672 13526 2688
rect 13909 3180 13963 3196
rect 13909 3146 13929 3180
rect 13909 3097 13963 3146
rect 13909 3063 13929 3097
rect 13909 3014 13963 3063
rect 13909 2980 13929 3014
rect 14003 3180 14069 3249
rect 14003 3146 14019 3180
rect 14053 3146 14069 3180
rect 14508 3176 14574 3249
rect 14003 3112 14069 3146
rect 14003 3078 14019 3112
rect 14053 3078 14069 3112
rect 14003 3044 14069 3078
rect 14003 3010 14019 3044
rect 14053 3010 14069 3044
rect 14308 3135 14374 3151
rect 14308 3101 14324 3135
rect 14358 3101 14374 3135
rect 14308 3067 14374 3101
rect 14308 3033 14324 3067
rect 14358 3033 14374 3067
rect 14308 3024 14374 3033
rect 13909 2964 13963 2980
rect 14103 2999 14374 3024
rect 14103 2990 14324 2999
rect 14103 2976 14137 2990
rect 13909 2826 13943 2964
rect 13999 2942 14137 2976
rect 14308 2965 14324 2990
rect 14358 2965 14374 2999
rect 14414 3135 14464 3151
rect 14448 3101 14464 3135
rect 14508 3142 14524 3176
rect 14558 3142 14574 3176
rect 14508 3126 14574 3142
rect 14414 3092 14464 3101
rect 14612 3108 14678 3151
rect 14612 3092 14628 3108
rect 14414 3074 14628 3092
rect 14662 3074 14678 3108
rect 14414 3058 14678 3074
rect 14713 3111 14779 3249
rect 14713 3077 14729 3111
rect 14763 3077 14779 3111
rect 14713 3061 14779 3077
rect 14906 3135 14991 3151
rect 14906 3101 14922 3135
rect 14956 3101 14991 3135
rect 14414 3043 14464 3058
rect 14448 3009 14464 3043
rect 14906 3024 14991 3101
rect 14414 2993 14464 3009
rect 14205 2950 14251 2956
rect 13999 2926 14033 2942
rect 13977 2910 14033 2926
rect 14011 2876 14033 2910
rect 14205 2916 14211 2950
rect 14245 2916 14251 2950
rect 14308 2949 14374 2965
rect 14498 2990 14922 3024
rect 14956 2990 14991 3024
rect 15025 3135 15082 3151
rect 15025 3101 15041 3135
rect 15075 3101 15082 3135
rect 15025 3051 15082 3101
rect 15116 3137 15257 3249
rect 15443 3180 15509 3249
rect 15954 3245 15985 3279
rect 16019 3245 16081 3279
rect 16115 3245 16177 3279
rect 16211 3245 16273 3279
rect 16307 3245 16369 3279
rect 16403 3245 16465 3279
rect 16499 3245 16561 3279
rect 16595 3245 16657 3279
rect 16691 3245 16753 3279
rect 16787 3245 16849 3279
rect 16883 3245 16945 3279
rect 16979 3245 17041 3279
rect 17075 3245 17137 3279
rect 17171 3245 17233 3279
rect 17267 3245 17329 3279
rect 17363 3245 17425 3279
rect 17459 3245 17521 3279
rect 17555 3245 17617 3279
rect 17651 3245 17682 3279
rect 15116 3103 15132 3137
rect 15166 3103 15207 3137
rect 15241 3103 15257 3137
rect 15116 3100 15257 3103
rect 15292 3150 15356 3166
rect 15292 3116 15306 3150
rect 15340 3116 15356 3150
rect 15292 3051 15356 3116
rect 15025 3017 15041 3051
rect 15075 3040 15356 3051
rect 15075 3017 15306 3040
rect 15290 3006 15306 3017
rect 15340 3006 15356 3040
rect 15290 2990 15356 3006
rect 15443 3146 15459 3180
rect 15493 3146 15509 3180
rect 15443 3097 15509 3146
rect 15443 3063 15459 3097
rect 15493 3063 15509 3097
rect 15443 3014 15509 3063
rect 14498 2959 14532 2990
rect 14205 2915 14251 2916
rect 14408 2925 14532 2959
rect 14957 2983 14991 2990
rect 14660 2950 14731 2956
rect 14408 2915 14442 2925
rect 13977 2860 14033 2876
rect 13909 2810 13965 2826
rect 13909 2776 13931 2810
rect 13909 2720 13965 2776
rect 13909 2686 13931 2720
rect 13999 2750 14033 2860
rect 14069 2894 14135 2908
rect 14069 2860 14085 2894
rect 14119 2860 14135 2894
rect 14069 2844 14135 2860
rect 14205 2899 14315 2915
rect 14205 2865 14265 2899
rect 14299 2865 14315 2899
rect 14205 2852 14315 2865
rect 14357 2899 14442 2915
rect 14357 2865 14373 2899
rect 14407 2865 14442 2899
rect 14660 2916 14691 2950
rect 14725 2916 14731 2950
rect 14660 2899 14731 2916
rect 14357 2852 14442 2865
rect 14552 2875 14618 2891
rect 14101 2818 14135 2844
rect 14552 2841 14568 2875
rect 14602 2841 14618 2875
rect 14660 2865 14676 2899
rect 14710 2865 14731 2899
rect 14877 2950 14923 2956
rect 14877 2916 14883 2950
rect 14917 2916 14923 2950
rect 14957 2949 15202 2983
rect 15443 2980 15459 3014
rect 15493 2980 15509 3014
rect 15443 2964 15509 2980
rect 15549 3180 15600 3196
rect 15583 3146 15600 3180
rect 15549 3097 15600 3146
rect 15583 3063 15600 3097
rect 15549 3014 15600 3063
rect 15583 2980 15600 3014
rect 14877 2915 14923 2916
rect 14877 2899 15020 2915
rect 14660 2852 14731 2865
rect 14768 2876 14834 2891
rect 14768 2875 14790 2876
rect 14552 2818 14618 2841
rect 14768 2841 14784 2875
rect 14824 2842 14834 2876
rect 14877 2865 14970 2899
rect 15004 2865 15020 2899
rect 14877 2855 15020 2865
rect 15054 2899 15134 2915
rect 15054 2865 15084 2899
rect 15118 2865 15134 2899
rect 15054 2864 15134 2865
rect 14818 2841 14834 2842
rect 14768 2821 14834 2841
rect 15054 2821 15088 2864
rect 15168 2830 15202 2949
rect 15252 2920 15386 2956
rect 15252 2914 15314 2920
rect 15354 2914 15386 2920
rect 15252 2880 15268 2914
rect 15302 2880 15314 2914
rect 15370 2880 15386 2914
rect 15549 2940 15600 2980
rect 15971 3176 16025 3192
rect 15971 3142 15991 3176
rect 15971 3093 16025 3142
rect 15971 3059 15991 3093
rect 15971 3010 16025 3059
rect 15971 2976 15991 3010
rect 16065 3176 16131 3245
rect 16065 3142 16081 3176
rect 16115 3142 16131 3176
rect 16570 3172 16636 3245
rect 16065 3108 16131 3142
rect 16065 3074 16081 3108
rect 16115 3074 16131 3108
rect 16065 3040 16131 3074
rect 16065 3006 16081 3040
rect 16115 3006 16131 3040
rect 16370 3131 16436 3147
rect 16370 3097 16386 3131
rect 16420 3097 16436 3131
rect 16370 3063 16436 3097
rect 16370 3029 16386 3063
rect 16420 3029 16436 3063
rect 16370 3020 16436 3029
rect 15971 2960 16025 2976
rect 16165 2995 16436 3020
rect 16165 2986 16386 2995
rect 16165 2972 16199 2986
rect 15252 2878 15314 2880
rect 15354 2878 15386 2880
rect 15252 2864 15386 2878
rect 15434 2894 15500 2910
rect 15434 2860 15450 2894
rect 15484 2860 15500 2894
rect 15434 2830 15500 2860
rect 14768 2818 15088 2821
rect 14101 2787 15088 2818
rect 15122 2796 15500 2830
rect 15549 2906 15568 2940
rect 15549 2826 15600 2906
rect 15534 2810 15600 2826
rect 14101 2784 14834 2787
rect 15122 2753 15156 2796
rect 15534 2776 15550 2810
rect 15584 2776 15600 2810
rect 13999 2727 14346 2750
rect 13999 2716 14296 2727
rect 13909 2670 13965 2686
rect 14280 2693 14296 2716
rect 14330 2693 14346 2727
rect 14017 2648 14035 2682
rect 14069 2648 14088 2682
rect 14280 2671 14346 2693
rect 14388 2734 14674 2750
rect 14388 2700 14412 2734
rect 14446 2716 14624 2734
rect 14446 2700 14470 2716
rect 14388 2684 14470 2700
rect 14608 2700 14624 2716
rect 14658 2700 14674 2734
rect 14608 2684 14674 2700
rect 14708 2726 14803 2742
rect 14708 2692 14738 2726
rect 14772 2692 14803 2726
rect 11818 2585 11849 2619
rect 11883 2585 11945 2619
rect 11979 2585 12041 2619
rect 12075 2585 12137 2619
rect 12171 2585 12233 2619
rect 12267 2585 12329 2619
rect 12363 2585 12425 2619
rect 12459 2585 12521 2619
rect 12555 2585 12617 2619
rect 12651 2585 12713 2619
rect 12747 2585 12809 2619
rect 12843 2585 12905 2619
rect 12939 2585 13001 2619
rect 13035 2585 13097 2619
rect 13131 2585 13193 2619
rect 13227 2585 13289 2619
rect 13323 2585 13385 2619
rect 13419 2585 13481 2619
rect 13515 2585 13546 2619
rect 14017 2617 14088 2648
rect 14506 2648 14522 2682
rect 14556 2648 14572 2682
rect 14506 2617 14572 2648
rect 14708 2617 14803 2692
rect 14901 2737 15156 2753
rect 14901 2703 14917 2737
rect 14951 2719 15156 2737
rect 15190 2746 15410 2762
rect 15190 2728 15360 2746
rect 14951 2703 14967 2719
rect 14901 2687 14967 2703
rect 15190 2685 15224 2728
rect 15344 2712 15360 2728
rect 15394 2712 15410 2746
rect 15344 2696 15410 2712
rect 15448 2738 15498 2754
rect 15448 2704 15464 2738
rect 15003 2651 15019 2685
rect 15053 2651 15113 2685
rect 15147 2651 15224 2685
rect 15258 2678 15308 2694
rect 15292 2644 15308 2678
rect 15258 2617 15308 2644
rect 15448 2617 15498 2704
rect 15534 2720 15600 2776
rect 15534 2686 15550 2720
rect 15584 2686 15600 2720
rect 15534 2670 15600 2686
rect 15971 2822 16005 2960
rect 16061 2938 16199 2972
rect 16370 2961 16386 2986
rect 16420 2961 16436 2995
rect 16476 3131 16526 3147
rect 16510 3097 16526 3131
rect 16570 3138 16586 3172
rect 16620 3138 16636 3172
rect 16570 3122 16636 3138
rect 16476 3088 16526 3097
rect 16674 3104 16740 3147
rect 16674 3088 16690 3104
rect 16476 3070 16690 3088
rect 16724 3070 16740 3104
rect 16476 3054 16740 3070
rect 16775 3107 16841 3245
rect 16775 3073 16791 3107
rect 16825 3073 16841 3107
rect 16775 3057 16841 3073
rect 16968 3131 17053 3147
rect 16968 3097 16984 3131
rect 17018 3097 17053 3131
rect 16476 3039 16526 3054
rect 16510 3005 16526 3039
rect 16968 3020 17053 3097
rect 16476 2989 16526 3005
rect 16267 2946 16313 2952
rect 16061 2922 16095 2938
rect 16039 2906 16095 2922
rect 16073 2872 16095 2906
rect 16267 2912 16273 2946
rect 16307 2912 16313 2946
rect 16370 2945 16436 2961
rect 16560 2986 16984 3020
rect 17018 2986 17053 3020
rect 17087 3131 17144 3147
rect 17087 3097 17103 3131
rect 17137 3097 17144 3131
rect 17087 3047 17144 3097
rect 17178 3133 17319 3245
rect 17505 3176 17571 3245
rect 17178 3099 17194 3133
rect 17228 3099 17269 3133
rect 17303 3099 17319 3133
rect 17178 3096 17319 3099
rect 17354 3146 17418 3162
rect 17354 3112 17368 3146
rect 17402 3112 17418 3146
rect 17354 3047 17418 3112
rect 17087 3013 17103 3047
rect 17137 3036 17418 3047
rect 17137 3013 17368 3036
rect 17352 3002 17368 3013
rect 17402 3002 17418 3036
rect 17352 2986 17418 3002
rect 17505 3142 17521 3176
rect 17555 3142 17571 3176
rect 17505 3093 17571 3142
rect 17505 3059 17521 3093
rect 17555 3059 17571 3093
rect 17505 3010 17571 3059
rect 16560 2955 16594 2986
rect 16267 2911 16313 2912
rect 16470 2921 16594 2955
rect 17019 2979 17053 2986
rect 16722 2946 16793 2952
rect 16470 2911 16504 2921
rect 16039 2856 16095 2872
rect 15971 2806 16027 2822
rect 15971 2772 15993 2806
rect 15971 2716 16027 2772
rect 15971 2682 15993 2716
rect 16061 2746 16095 2856
rect 16131 2890 16197 2904
rect 16131 2856 16147 2890
rect 16181 2856 16197 2890
rect 16131 2840 16197 2856
rect 16267 2895 16377 2911
rect 16267 2861 16327 2895
rect 16361 2861 16377 2895
rect 16267 2848 16377 2861
rect 16419 2895 16504 2911
rect 16419 2861 16435 2895
rect 16469 2861 16504 2895
rect 16722 2912 16753 2946
rect 16787 2912 16793 2946
rect 16722 2895 16793 2912
rect 16419 2848 16504 2861
rect 16614 2871 16680 2887
rect 16163 2814 16197 2840
rect 16614 2837 16630 2871
rect 16664 2837 16680 2871
rect 16722 2861 16738 2895
rect 16772 2861 16793 2895
rect 16939 2946 16985 2952
rect 16939 2912 16945 2946
rect 16979 2912 16985 2946
rect 17019 2945 17264 2979
rect 17505 2976 17521 3010
rect 17555 2976 17571 3010
rect 17505 2960 17571 2976
rect 17611 3176 17662 3192
rect 17645 3142 17662 3176
rect 17611 3093 17662 3142
rect 17645 3059 17662 3093
rect 17611 3010 17662 3059
rect 17645 2976 17662 3010
rect 16939 2911 16985 2912
rect 16939 2895 17082 2911
rect 16722 2848 16793 2861
rect 16830 2872 16896 2887
rect 16830 2871 16852 2872
rect 16614 2814 16680 2837
rect 16830 2837 16846 2871
rect 16886 2838 16896 2872
rect 16939 2861 17032 2895
rect 17066 2861 17082 2895
rect 16939 2851 17082 2861
rect 17116 2895 17196 2911
rect 17116 2861 17146 2895
rect 17180 2861 17196 2895
rect 17116 2860 17196 2861
rect 16880 2837 16896 2838
rect 16830 2817 16896 2837
rect 17116 2817 17150 2860
rect 17230 2826 17264 2945
rect 17314 2916 17448 2952
rect 17314 2910 17376 2916
rect 17416 2910 17448 2916
rect 17314 2876 17330 2910
rect 17364 2876 17376 2910
rect 17432 2876 17448 2910
rect 17314 2874 17376 2876
rect 17416 2874 17448 2876
rect 17314 2860 17448 2874
rect 17496 2890 17562 2906
rect 17496 2856 17512 2890
rect 17546 2856 17562 2890
rect 17496 2826 17562 2856
rect 16830 2814 17150 2817
rect 16163 2783 17150 2814
rect 17184 2792 17562 2826
rect 17611 2846 17662 2976
rect 17611 2822 17616 2846
rect 17596 2808 17616 2822
rect 17658 2808 17662 2846
rect 17596 2806 17662 2808
rect 16163 2780 16896 2783
rect 17184 2749 17218 2792
rect 17596 2772 17612 2806
rect 17646 2772 17662 2806
rect 16061 2723 16408 2746
rect 16061 2712 16358 2723
rect 15971 2666 16027 2682
rect 16342 2689 16358 2712
rect 16392 2689 16408 2723
rect 16079 2644 16097 2678
rect 16131 2644 16150 2678
rect 16342 2667 16408 2689
rect 16450 2730 16736 2746
rect 16450 2696 16474 2730
rect 16508 2712 16686 2730
rect 16508 2696 16532 2712
rect 16450 2680 16532 2696
rect 16670 2696 16686 2712
rect 16720 2696 16736 2730
rect 16670 2680 16736 2696
rect 16770 2722 16865 2738
rect 16770 2688 16800 2722
rect 16834 2688 16865 2722
rect 13892 2583 13923 2617
rect 13957 2583 14019 2617
rect 14053 2583 14115 2617
rect 14149 2583 14211 2617
rect 14245 2583 14307 2617
rect 14341 2583 14403 2617
rect 14437 2583 14499 2617
rect 14533 2583 14595 2617
rect 14629 2583 14691 2617
rect 14725 2583 14787 2617
rect 14821 2583 14883 2617
rect 14917 2583 14979 2617
rect 15013 2583 15075 2617
rect 15109 2583 15171 2617
rect 15205 2583 15267 2617
rect 15301 2583 15363 2617
rect 15397 2583 15459 2617
rect 15493 2583 15555 2617
rect 15589 2583 15620 2617
rect 16079 2613 16150 2644
rect 16568 2644 16584 2678
rect 16618 2644 16634 2678
rect 16568 2613 16634 2644
rect 16770 2613 16865 2688
rect 16963 2733 17218 2749
rect 16963 2699 16979 2733
rect 17013 2715 17218 2733
rect 17252 2742 17472 2758
rect 17252 2724 17422 2742
rect 17013 2699 17029 2715
rect 16963 2683 17029 2699
rect 17252 2681 17286 2724
rect 17406 2708 17422 2724
rect 17456 2708 17472 2742
rect 17406 2692 17472 2708
rect 17510 2734 17560 2750
rect 17510 2700 17526 2734
rect 17065 2647 17081 2681
rect 17115 2647 17175 2681
rect 17209 2647 17286 2681
rect 17320 2674 17370 2690
rect 17354 2640 17370 2674
rect 17320 2613 17370 2640
rect 17510 2613 17560 2700
rect 17596 2716 17662 2772
rect 17596 2682 17612 2716
rect 17646 2682 17662 2716
rect 17596 2666 17662 2682
rect 15954 2579 15985 2613
rect 16019 2579 16081 2613
rect 16115 2579 16177 2613
rect 16211 2579 16273 2613
rect 16307 2579 16369 2613
rect 16403 2579 16465 2613
rect 16499 2579 16561 2613
rect 16595 2579 16657 2613
rect 16691 2579 16753 2613
rect 16787 2579 16849 2613
rect 16883 2579 16945 2613
rect 16979 2579 17041 2613
rect 17075 2579 17137 2613
rect 17171 2579 17233 2613
rect 17267 2579 17329 2613
rect 17363 2579 17425 2613
rect 17459 2579 17521 2613
rect 17555 2579 17617 2613
rect 17651 2579 17682 2613
<< viali >>
rect 18151 6127 18185 6161
rect 18243 6127 18277 6161
rect 18335 6127 18369 6161
rect 26321 6079 26355 6113
rect 26413 6079 26447 6113
rect 26505 6079 26539 6113
rect 26597 6079 26631 6113
rect 26689 6079 26723 6113
rect 26781 6079 26815 6113
rect 26873 6079 26907 6113
rect 26965 6079 26999 6113
rect 27057 6079 27091 6113
rect 27149 6079 27183 6113
rect 27241 6079 27275 6113
rect 27333 6079 27367 6113
rect 27425 6079 27459 6113
rect 27517 6079 27551 6113
rect 27609 6079 27643 6113
rect 27701 6079 27735 6113
rect 18196 5849 18236 5854
rect 18196 5816 18202 5849
rect 18202 5816 18236 5849
rect 18298 5818 18332 5852
rect 28127 6061 28161 6095
rect 28219 6061 28253 6095
rect 28311 6061 28345 6095
rect 28403 6061 28437 6095
rect 28495 6061 28529 6095
rect 28587 6061 28621 6095
rect 28679 6061 28713 6095
rect 28771 6061 28805 6095
rect 28863 6061 28897 6095
rect 28955 6061 28989 6095
rect 29047 6061 29081 6095
rect 29139 6061 29173 6095
rect 29231 6061 29265 6095
rect 29323 6061 29357 6095
rect 29415 6061 29449 6095
rect 29507 6061 29541 6095
rect 17028 5742 17068 5778
rect 18818 5802 18858 5840
rect 18920 5804 18954 5838
rect 19396 5804 19430 5838
rect 19498 5790 19532 5824
rect 20032 5788 20066 5822
rect 20374 5784 20408 5818
rect 17302 5700 17354 5752
rect 17416 5696 17468 5748
rect 20842 5776 20882 5814
rect 21382 5780 21418 5820
rect 21954 5782 21992 5824
rect 22548 5776 22590 5818
rect 23136 5782 23174 5824
rect 24080 5768 24122 5806
rect 24520 5766 24562 5804
rect 25776 5766 25818 5804
rect 26364 5801 26406 5810
rect 26364 5772 26368 5801
rect 26368 5772 26406 5801
rect 27600 5756 27640 5794
rect 28170 5783 28212 5792
rect 28170 5754 28174 5783
rect 28174 5754 28212 5783
rect 18151 5583 18185 5617
rect 18243 5583 18277 5617
rect 18335 5583 18369 5617
rect 29406 5738 29446 5776
rect 26321 5535 26355 5569
rect 26413 5535 26447 5569
rect 26505 5535 26539 5569
rect 26597 5535 26631 5569
rect 26689 5535 26723 5569
rect 26781 5535 26815 5569
rect 26873 5535 26907 5569
rect 26965 5535 26999 5569
rect 27057 5535 27091 5569
rect 27149 5535 27183 5569
rect 27241 5535 27275 5569
rect 27333 5535 27367 5569
rect 27425 5535 27459 5569
rect 27517 5535 27551 5569
rect 27609 5535 27643 5569
rect 27701 5535 27735 5569
rect 28127 5517 28161 5551
rect 28219 5517 28253 5551
rect 28311 5517 28345 5551
rect 28403 5517 28437 5551
rect 28495 5517 28529 5551
rect 28587 5517 28621 5551
rect 28679 5517 28713 5551
rect 28771 5517 28805 5551
rect 28863 5517 28897 5551
rect 28955 5517 28989 5551
rect 29047 5517 29081 5551
rect 29139 5517 29173 5551
rect 29231 5517 29265 5551
rect 29323 5517 29357 5551
rect 29415 5517 29449 5551
rect 29507 5517 29541 5551
rect 8220 4096 8256 4138
rect 8320 4112 8354 4146
rect 1529 3269 1563 3303
rect 1625 3269 1659 3303
rect 1721 3269 1755 3303
rect 1817 3269 1851 3303
rect 1913 3269 1947 3303
rect 2009 3269 2043 3303
rect 2105 3269 2139 3303
rect 2201 3269 2235 3303
rect 2297 3269 2331 3303
rect 2393 3269 2427 3303
rect 2489 3269 2523 3303
rect 2585 3269 2619 3303
rect 2681 3269 2715 3303
rect 2777 3269 2811 3303
rect 2873 3269 2907 3303
rect 2969 3269 3003 3303
rect 3065 3269 3099 3303
rect 3161 3269 3195 3303
rect 1817 2936 1851 2970
rect 3591 3265 3625 3299
rect 3687 3265 3721 3299
rect 3783 3265 3817 3299
rect 3879 3265 3913 3299
rect 3975 3265 4009 3299
rect 4071 3265 4105 3299
rect 4167 3265 4201 3299
rect 4263 3265 4297 3299
rect 4359 3265 4393 3299
rect 4455 3265 4489 3299
rect 4551 3265 4585 3299
rect 4647 3265 4681 3299
rect 4743 3265 4777 3299
rect 4839 3265 4873 3299
rect 4935 3265 4969 3299
rect 5031 3265 5065 3299
rect 5127 3265 5161 3299
rect 5223 3265 5257 3299
rect 2297 2936 2331 2970
rect 2489 2936 2523 2970
rect 2396 2895 2430 2896
rect 2396 2862 2424 2895
rect 2424 2862 2430 2895
rect 2920 2934 2960 2940
rect 2920 2900 2942 2934
rect 2942 2900 2960 2934
rect 2920 2898 2960 2900
rect 3174 2926 3208 2960
rect 3879 2932 3913 2966
rect 5665 3263 5699 3297
rect 5761 3263 5795 3297
rect 5857 3263 5891 3297
rect 5953 3263 5987 3297
rect 6049 3263 6083 3297
rect 6145 3263 6179 3297
rect 6241 3263 6275 3297
rect 6337 3263 6371 3297
rect 6433 3263 6467 3297
rect 6529 3263 6563 3297
rect 6625 3263 6659 3297
rect 6721 3263 6755 3297
rect 6817 3263 6851 3297
rect 6913 3263 6947 3297
rect 7009 3263 7043 3297
rect 7105 3263 7139 3297
rect 7201 3263 7235 3297
rect 7297 3263 7331 3297
rect 4359 2932 4393 2966
rect 4551 2932 4585 2966
rect 4458 2891 4492 2892
rect 4458 2858 4486 2891
rect 4486 2858 4492 2891
rect 4982 2930 5022 2936
rect 4982 2896 5004 2930
rect 5004 2896 5022 2930
rect 5232 2928 5268 2962
rect 4982 2894 5022 2896
rect 1529 2603 1563 2637
rect 1625 2603 1659 2637
rect 1721 2603 1755 2637
rect 1817 2603 1851 2637
rect 1913 2603 1947 2637
rect 2009 2603 2043 2637
rect 2105 2603 2139 2637
rect 2201 2603 2235 2637
rect 2297 2603 2331 2637
rect 2393 2603 2427 2637
rect 2489 2603 2523 2637
rect 2585 2603 2619 2637
rect 2681 2603 2715 2637
rect 2777 2603 2811 2637
rect 2873 2603 2907 2637
rect 2969 2603 3003 2637
rect 3065 2603 3099 2637
rect 3161 2603 3195 2637
rect 5953 2930 5987 2964
rect 7727 3259 7761 3293
rect 7823 3259 7857 3293
rect 7919 3259 7953 3293
rect 8015 3259 8049 3293
rect 8111 3259 8145 3293
rect 8207 3259 8241 3293
rect 8303 3259 8337 3293
rect 8399 3259 8433 3293
rect 8495 3259 8529 3293
rect 8591 3259 8625 3293
rect 8687 3259 8721 3293
rect 8783 3259 8817 3293
rect 8879 3259 8913 3293
rect 8975 3259 9009 3293
rect 9071 3259 9105 3293
rect 9167 3259 9201 3293
rect 9263 3259 9297 3293
rect 9359 3259 9393 3293
rect 6433 2930 6467 2964
rect 6625 2930 6659 2964
rect 6532 2889 6566 2890
rect 6532 2856 6560 2889
rect 6560 2856 6566 2889
rect 7056 2928 7096 2934
rect 7056 2894 7078 2928
rect 7078 2894 7096 2928
rect 7056 2892 7096 2894
rect 7310 2920 7344 2954
rect 3591 2599 3625 2633
rect 3687 2599 3721 2633
rect 3783 2599 3817 2633
rect 3879 2599 3913 2633
rect 3975 2599 4009 2633
rect 4071 2599 4105 2633
rect 4167 2599 4201 2633
rect 4263 2599 4297 2633
rect 4359 2599 4393 2633
rect 4455 2599 4489 2633
rect 4551 2599 4585 2633
rect 4647 2599 4681 2633
rect 4743 2599 4777 2633
rect 4839 2599 4873 2633
rect 4935 2599 4969 2633
rect 5031 2599 5065 2633
rect 5127 2599 5161 2633
rect 5223 2599 5257 2633
rect 8015 2926 8049 2960
rect 9787 3255 9821 3289
rect 9883 3255 9917 3289
rect 9979 3255 10013 3289
rect 10075 3255 10109 3289
rect 10171 3255 10205 3289
rect 10267 3255 10301 3289
rect 10363 3255 10397 3289
rect 10459 3255 10493 3289
rect 10555 3255 10589 3289
rect 10651 3255 10685 3289
rect 10747 3255 10781 3289
rect 10843 3255 10877 3289
rect 10939 3255 10973 3289
rect 11035 3255 11069 3289
rect 11131 3255 11165 3289
rect 11227 3255 11261 3289
rect 11323 3255 11357 3289
rect 11419 3255 11453 3289
rect 8495 2926 8529 2960
rect 8687 2926 8721 2960
rect 8594 2885 8628 2886
rect 8594 2852 8622 2885
rect 8622 2852 8628 2885
rect 9118 2924 9158 2930
rect 9118 2890 9140 2924
rect 9140 2890 9158 2924
rect 9118 2888 9158 2890
rect 9366 2910 9402 2944
rect 5665 2597 5699 2631
rect 5761 2597 5795 2631
rect 5857 2597 5891 2631
rect 5953 2597 5987 2631
rect 6049 2597 6083 2631
rect 6145 2597 6179 2631
rect 6241 2597 6275 2631
rect 6337 2597 6371 2631
rect 6433 2597 6467 2631
rect 6529 2597 6563 2631
rect 6625 2597 6659 2631
rect 6721 2597 6755 2631
rect 6817 2597 6851 2631
rect 6913 2597 6947 2631
rect 7009 2597 7043 2631
rect 7105 2597 7139 2631
rect 7201 2597 7235 2631
rect 7297 2597 7331 2631
rect 10075 2922 10109 2956
rect 11849 3251 11883 3285
rect 11945 3251 11979 3285
rect 12041 3251 12075 3285
rect 12137 3251 12171 3285
rect 12233 3251 12267 3285
rect 12329 3251 12363 3285
rect 12425 3251 12459 3285
rect 12521 3251 12555 3285
rect 12617 3251 12651 3285
rect 12713 3251 12747 3285
rect 12809 3251 12843 3285
rect 12905 3251 12939 3285
rect 13001 3251 13035 3285
rect 13097 3251 13131 3285
rect 13193 3251 13227 3285
rect 13289 3251 13323 3285
rect 13385 3251 13419 3285
rect 13481 3251 13515 3285
rect 10555 2922 10589 2956
rect 10747 2922 10781 2956
rect 10654 2881 10688 2882
rect 10654 2848 10682 2881
rect 10682 2848 10688 2881
rect 11178 2920 11218 2926
rect 11178 2886 11200 2920
rect 11200 2886 11218 2920
rect 11178 2884 11218 2886
rect 11432 2912 11466 2946
rect 7727 2593 7761 2627
rect 7823 2593 7857 2627
rect 7919 2593 7953 2627
rect 8015 2593 8049 2627
rect 8111 2593 8145 2627
rect 8207 2593 8241 2627
rect 8303 2593 8337 2627
rect 8399 2593 8433 2627
rect 8495 2593 8529 2627
rect 8591 2593 8625 2627
rect 8687 2593 8721 2627
rect 8783 2593 8817 2627
rect 8879 2593 8913 2627
rect 8975 2593 9009 2627
rect 9071 2593 9105 2627
rect 9167 2593 9201 2627
rect 9263 2593 9297 2627
rect 9359 2593 9393 2627
rect 12137 2918 12171 2952
rect 13923 3249 13957 3283
rect 14019 3249 14053 3283
rect 14115 3249 14149 3283
rect 14211 3249 14245 3283
rect 14307 3249 14341 3283
rect 14403 3249 14437 3283
rect 14499 3249 14533 3283
rect 14595 3249 14629 3283
rect 14691 3249 14725 3283
rect 14787 3249 14821 3283
rect 14883 3249 14917 3283
rect 14979 3249 15013 3283
rect 15075 3249 15109 3283
rect 15171 3249 15205 3283
rect 15267 3249 15301 3283
rect 15363 3249 15397 3283
rect 15459 3249 15493 3283
rect 15555 3249 15589 3283
rect 12617 2918 12651 2952
rect 12809 2918 12843 2952
rect 12716 2877 12750 2878
rect 12716 2844 12744 2877
rect 12744 2844 12750 2877
rect 13240 2916 13280 2922
rect 13240 2882 13262 2916
rect 13262 2882 13280 2916
rect 13490 2914 13526 2948
rect 13240 2880 13280 2882
rect 9787 2589 9821 2623
rect 9883 2589 9917 2623
rect 9979 2589 10013 2623
rect 10075 2589 10109 2623
rect 10171 2589 10205 2623
rect 10267 2589 10301 2623
rect 10363 2589 10397 2623
rect 10459 2589 10493 2623
rect 10555 2589 10589 2623
rect 10651 2589 10685 2623
rect 10747 2589 10781 2623
rect 10843 2589 10877 2623
rect 10939 2589 10973 2623
rect 11035 2589 11069 2623
rect 11131 2589 11165 2623
rect 11227 2589 11261 2623
rect 11323 2589 11357 2623
rect 11419 2589 11453 2623
rect 14211 2916 14245 2950
rect 15985 3245 16019 3279
rect 16081 3245 16115 3279
rect 16177 3245 16211 3279
rect 16273 3245 16307 3279
rect 16369 3245 16403 3279
rect 16465 3245 16499 3279
rect 16561 3245 16595 3279
rect 16657 3245 16691 3279
rect 16753 3245 16787 3279
rect 16849 3245 16883 3279
rect 16945 3245 16979 3279
rect 17041 3245 17075 3279
rect 17137 3245 17171 3279
rect 17233 3245 17267 3279
rect 17329 3245 17363 3279
rect 17425 3245 17459 3279
rect 17521 3245 17555 3279
rect 17617 3245 17651 3279
rect 14691 2916 14725 2950
rect 14883 2916 14917 2950
rect 14790 2875 14824 2876
rect 14790 2842 14818 2875
rect 14818 2842 14824 2875
rect 15314 2914 15354 2920
rect 15314 2880 15336 2914
rect 15336 2880 15354 2914
rect 15314 2878 15354 2880
rect 15568 2906 15602 2940
rect 11849 2585 11883 2619
rect 11945 2585 11979 2619
rect 12041 2585 12075 2619
rect 12137 2585 12171 2619
rect 12233 2585 12267 2619
rect 12329 2585 12363 2619
rect 12425 2585 12459 2619
rect 12521 2585 12555 2619
rect 12617 2585 12651 2619
rect 12713 2585 12747 2619
rect 12809 2585 12843 2619
rect 12905 2585 12939 2619
rect 13001 2585 13035 2619
rect 13097 2585 13131 2619
rect 13193 2585 13227 2619
rect 13289 2585 13323 2619
rect 13385 2585 13419 2619
rect 13481 2585 13515 2619
rect 16273 2912 16307 2946
rect 16753 2912 16787 2946
rect 16945 2912 16979 2946
rect 16852 2871 16886 2872
rect 16852 2838 16880 2871
rect 16880 2838 16886 2871
rect 17376 2910 17416 2916
rect 17376 2876 17398 2910
rect 17398 2876 17416 2910
rect 17376 2874 17416 2876
rect 17616 2808 17658 2846
rect 13923 2583 13957 2617
rect 14019 2583 14053 2617
rect 14115 2583 14149 2617
rect 14211 2583 14245 2617
rect 14307 2583 14341 2617
rect 14403 2583 14437 2617
rect 14499 2583 14533 2617
rect 14595 2583 14629 2617
rect 14691 2583 14725 2617
rect 14787 2583 14821 2617
rect 14883 2583 14917 2617
rect 14979 2583 15013 2617
rect 15075 2583 15109 2617
rect 15171 2583 15205 2617
rect 15267 2583 15301 2617
rect 15363 2583 15397 2617
rect 15459 2583 15493 2617
rect 15555 2583 15589 2617
rect 15985 2579 16019 2613
rect 16081 2579 16115 2613
rect 16177 2579 16211 2613
rect 16273 2579 16307 2613
rect 16369 2579 16403 2613
rect 16465 2579 16499 2613
rect 16561 2579 16595 2613
rect 16657 2579 16691 2613
rect 16753 2579 16787 2613
rect 16849 2579 16883 2613
rect 16945 2579 16979 2613
rect 17041 2579 17075 2613
rect 17137 2579 17171 2613
rect 17233 2579 17267 2613
rect 17329 2579 17363 2613
rect 17425 2579 17459 2613
rect 17521 2579 17555 2613
rect 17617 2579 17651 2613
<< metal1 >>
rect 27624 45014 27752 45042
rect 27624 44952 27662 45014
rect 27722 44952 27752 45014
rect 27624 44946 27752 44952
rect 27624 9475 27662 44946
rect 16465 9437 27662 9475
rect 16465 5763 16503 9437
rect 18122 6172 18398 6192
rect 18122 6161 18232 6172
rect 18284 6161 18398 6172
rect 18122 6127 18151 6161
rect 18185 6127 18232 6161
rect 18284 6127 18335 6161
rect 18369 6127 18398 6161
rect 18122 6120 18232 6127
rect 18284 6120 18398 6127
rect 18122 6096 18398 6120
rect 26292 6113 27032 6144
rect 27086 6113 27764 6144
rect 26292 6079 26321 6113
rect 26355 6079 26413 6113
rect 26447 6079 26505 6113
rect 26539 6079 26597 6113
rect 26631 6079 26689 6113
rect 26723 6079 26781 6113
rect 26815 6079 26873 6113
rect 26907 6079 26965 6113
rect 26999 6092 27032 6113
rect 26999 6079 27057 6092
rect 27091 6079 27149 6113
rect 27183 6079 27241 6113
rect 27275 6079 27333 6113
rect 27367 6079 27425 6113
rect 27459 6079 27517 6113
rect 27551 6079 27609 6113
rect 27643 6079 27701 6113
rect 27735 6079 27764 6113
rect 26292 6048 27764 6079
rect 28098 6095 28838 6126
rect 28892 6095 29570 6126
rect 28098 6061 28127 6095
rect 28161 6061 28219 6095
rect 28253 6061 28311 6095
rect 28345 6061 28403 6095
rect 28437 6061 28495 6095
rect 28529 6061 28587 6095
rect 28621 6061 28679 6095
rect 28713 6061 28771 6095
rect 28805 6074 28838 6095
rect 28805 6061 28863 6074
rect 28897 6061 28955 6095
rect 28989 6061 29047 6095
rect 29081 6061 29139 6095
rect 29173 6061 29231 6095
rect 29265 6061 29323 6095
rect 29357 6061 29415 6095
rect 29449 6061 29507 6095
rect 29541 6061 29570 6095
rect 28098 6030 29570 6061
rect 18064 5876 18450 5890
rect 18064 5860 20476 5876
rect 18064 5854 20516 5860
rect 18064 5816 18196 5854
rect 18236 5852 20516 5854
rect 18236 5818 18298 5852
rect 18332 5840 20516 5852
rect 18332 5818 18818 5840
rect 18236 5816 18818 5818
rect 18064 5802 18818 5816
rect 18858 5838 20516 5840
rect 18858 5804 18920 5838
rect 18954 5804 19396 5838
rect 19430 5824 20516 5838
rect 19430 5804 19498 5824
rect 18858 5802 19498 5804
rect 17019 5778 17088 5800
rect 17019 5763 17028 5778
rect 16465 5742 17028 5763
rect 17068 5742 17088 5778
rect 18064 5790 19498 5802
rect 19532 5822 20516 5824
rect 19532 5790 20032 5822
rect 18064 5788 20032 5790
rect 20066 5818 20516 5822
rect 20818 5818 20894 5846
rect 21371 5824 22057 5876
rect 21371 5820 21954 5824
rect 20066 5788 20374 5818
rect 18064 5784 20374 5788
rect 20408 5814 20918 5818
rect 20408 5784 20842 5814
rect 18064 5776 20842 5784
rect 20882 5776 20918 5814
rect 21371 5780 21382 5820
rect 21418 5782 21954 5820
rect 21992 5782 22057 5824
rect 21418 5780 22057 5782
rect 18064 5772 20476 5776
rect 16465 5730 17088 5742
rect 17292 5752 17374 5764
rect 16465 5725 17085 5730
rect 17292 5700 17302 5752
rect 17354 5700 17374 5752
rect 17292 5686 17374 5700
rect 17406 5748 17512 5760
rect 18388 5758 20476 5772
rect 20818 5756 20894 5776
rect 21371 5758 22057 5780
rect 22532 5824 23190 5832
rect 22532 5818 23136 5824
rect 22532 5776 22548 5818
rect 22590 5782 23136 5818
rect 23174 5782 23190 5824
rect 22590 5776 23190 5782
rect 22532 5766 23190 5776
rect 24068 5806 24634 5814
rect 24068 5768 24080 5806
rect 24122 5804 24634 5806
rect 24122 5768 24520 5804
rect 24068 5766 24520 5768
rect 24562 5766 24634 5804
rect 24068 5760 24634 5766
rect 25764 5810 26422 5822
rect 25764 5804 26364 5810
rect 25764 5766 25776 5804
rect 25818 5772 26364 5804
rect 26406 5772 26422 5810
rect 25818 5766 26422 5772
rect 25764 5754 26422 5766
rect 27590 5804 28009 5816
rect 27590 5794 28228 5804
rect 29608 5798 30506 5816
rect 27590 5756 27600 5794
rect 27640 5792 28228 5794
rect 27640 5756 28170 5792
rect 27590 5754 28170 5756
rect 28212 5754 28228 5792
rect 17406 5696 17416 5748
rect 17468 5696 17512 5748
rect 27590 5738 28228 5754
rect 27974 5736 28228 5738
rect 29396 5794 30506 5798
rect 29396 5776 30508 5794
rect 29396 5738 29406 5776
rect 29446 5738 30508 5776
rect 29396 5720 29614 5738
rect 17406 5670 17512 5696
rect 18122 5630 18398 5648
rect 18122 5617 18236 5630
rect 18290 5617 18398 5630
rect 18122 5583 18151 5617
rect 18185 5583 18236 5617
rect 18290 5583 18335 5617
rect 18369 5583 18398 5617
rect 18122 5570 18236 5583
rect 18290 5570 18398 5583
rect 18122 5552 18398 5570
rect 26292 5569 27764 5600
rect 26292 5535 26321 5569
rect 26355 5535 26413 5569
rect 26447 5535 26505 5569
rect 26539 5535 26597 5569
rect 26631 5535 26689 5569
rect 26723 5535 26781 5569
rect 26815 5535 26873 5569
rect 26907 5535 26965 5569
rect 26999 5564 27057 5569
rect 27091 5564 27149 5569
rect 26999 5535 27048 5564
rect 27104 5535 27149 5564
rect 27183 5535 27241 5569
rect 27275 5535 27333 5569
rect 27367 5535 27425 5569
rect 27459 5535 27517 5569
rect 27551 5535 27609 5569
rect 27643 5535 27701 5569
rect 27735 5535 27764 5569
rect 26292 5508 27048 5535
rect 27104 5508 27764 5535
rect 26292 5504 27764 5508
rect 28098 5551 29570 5582
rect 28098 5517 28127 5551
rect 28161 5517 28219 5551
rect 28253 5517 28311 5551
rect 28345 5517 28403 5551
rect 28437 5517 28495 5551
rect 28529 5517 28587 5551
rect 28621 5517 28679 5551
rect 28713 5517 28771 5551
rect 28805 5546 28863 5551
rect 28897 5546 28955 5551
rect 28805 5517 28854 5546
rect 28910 5517 28955 5546
rect 28989 5517 29047 5551
rect 29081 5517 29139 5551
rect 29173 5517 29231 5551
rect 29265 5517 29323 5551
rect 29357 5517 29415 5551
rect 29449 5517 29507 5551
rect 29541 5517 29570 5551
rect 28098 5490 28854 5517
rect 28910 5490 29570 5517
rect 28098 5486 29570 5490
rect 890 4486 972 4516
rect 890 4420 904 4486
rect 958 4473 972 4486
rect 958 4441 8130 4473
rect 958 4420 972 4441
rect 890 4386 972 4420
rect 8304 4196 8384 4204
rect 8182 4142 8266 4174
rect 8304 4158 8312 4196
rect 8182 4090 8192 4142
rect 8244 4138 8266 4142
rect 8256 4096 8266 4138
rect 8244 4090 8266 4096
rect 8182 4060 8266 4090
rect 8307 4144 8312 4158
rect 8364 4158 8384 4196
rect 8364 4144 8368 4158
rect 8307 4112 8320 4144
rect 8354 4112 8368 4144
rect 8307 4086 8368 4112
rect 8220 4044 8265 4060
rect 294 3830 484 3880
rect 294 3740 344 3830
rect 438 3807 484 3830
rect 438 3775 8130 3807
rect 438 3740 484 3775
rect 294 3684 484 3740
rect 1504 3332 3226 3335
rect 1504 3303 2482 3332
rect 2544 3308 3226 3332
rect 3560 3324 5288 3331
rect 3560 3308 4532 3324
rect 2544 3303 3232 3308
rect 1504 3269 1529 3303
rect 1563 3269 1625 3303
rect 1659 3269 1721 3303
rect 1755 3269 1817 3303
rect 1851 3269 1913 3303
rect 1947 3269 2009 3303
rect 2043 3269 2105 3303
rect 2139 3269 2201 3303
rect 2235 3269 2297 3303
rect 2331 3269 2393 3303
rect 2427 3270 2482 3303
rect 2544 3270 2585 3303
rect 2427 3269 2489 3270
rect 2523 3269 2585 3270
rect 2619 3269 2681 3303
rect 2715 3269 2777 3303
rect 2811 3269 2873 3303
rect 2907 3269 2969 3303
rect 3003 3269 3065 3303
rect 3099 3269 3161 3303
rect 3195 3269 3232 3303
rect 1504 3260 3232 3269
rect 3556 3299 4532 3308
rect 4594 3299 5288 3324
rect 3556 3265 3591 3299
rect 3625 3265 3687 3299
rect 3721 3265 3783 3299
rect 3817 3265 3879 3299
rect 3913 3265 3975 3299
rect 4009 3265 4071 3299
rect 4105 3265 4167 3299
rect 4201 3265 4263 3299
rect 4297 3265 4359 3299
rect 4393 3265 4455 3299
rect 4489 3265 4532 3299
rect 4594 3265 4647 3299
rect 4681 3265 4743 3299
rect 4777 3265 4839 3299
rect 4873 3265 4935 3299
rect 4969 3265 5031 3299
rect 5065 3265 5127 3299
rect 5161 3265 5223 3299
rect 5257 3298 5288 3299
rect 5634 3326 7362 3329
rect 5634 3298 6482 3326
rect 5257 3265 5292 3298
rect 3556 3262 4532 3265
rect 4594 3262 5292 3265
rect 3556 3260 5292 3262
rect 1504 3237 3226 3260
rect 3560 3250 5292 3260
rect 5616 3297 6482 3298
rect 6544 3298 7362 3326
rect 7696 3318 9424 3325
rect 7696 3298 8590 3318
rect 6544 3297 7364 3298
rect 5616 3263 5665 3297
rect 5699 3263 5761 3297
rect 5795 3263 5857 3297
rect 5891 3263 5953 3297
rect 5987 3263 6049 3297
rect 6083 3263 6145 3297
rect 6179 3263 6241 3297
rect 6275 3263 6337 3297
rect 6371 3263 6433 3297
rect 6467 3264 6482 3297
rect 6467 3263 6529 3264
rect 6563 3263 6625 3297
rect 6659 3263 6721 3297
rect 6755 3263 6817 3297
rect 6851 3263 6913 3297
rect 6947 3263 7009 3297
rect 7043 3263 7105 3297
rect 7139 3263 7201 3297
rect 7235 3263 7297 3297
rect 7331 3263 7364 3297
rect 5616 3250 7364 3263
rect 7688 3293 8590 3298
rect 8652 3293 9424 3318
rect 9756 3320 11484 3321
rect 9756 3300 10698 3320
rect 7688 3259 7727 3293
rect 7761 3259 7823 3293
rect 7857 3259 7919 3293
rect 7953 3259 8015 3293
rect 8049 3259 8111 3293
rect 8145 3259 8207 3293
rect 8241 3259 8303 3293
rect 8337 3259 8399 3293
rect 8433 3259 8495 3293
rect 8529 3259 8590 3293
rect 8652 3259 8687 3293
rect 8721 3259 8783 3293
rect 8817 3259 8879 3293
rect 8913 3259 8975 3293
rect 9009 3259 9071 3293
rect 9105 3259 9167 3293
rect 9201 3259 9263 3293
rect 9297 3259 9359 3293
rect 9393 3259 9424 3293
rect 7688 3256 8590 3259
rect 8652 3256 9424 3259
rect 7688 3250 9424 3256
rect 9748 3289 10698 3300
rect 10760 3289 11484 3320
rect 9748 3255 9787 3289
rect 9821 3255 9883 3289
rect 9917 3255 9979 3289
rect 10013 3255 10075 3289
rect 10109 3255 10171 3289
rect 10205 3255 10267 3289
rect 10301 3255 10363 3289
rect 10397 3255 10459 3289
rect 10493 3255 10555 3289
rect 10589 3255 10651 3289
rect 10685 3258 10698 3289
rect 10685 3255 10747 3258
rect 10781 3255 10843 3289
rect 10877 3255 10939 3289
rect 10973 3255 11035 3289
rect 11069 3255 11131 3289
rect 11165 3255 11227 3289
rect 11261 3255 11323 3289
rect 11357 3255 11419 3289
rect 11453 3286 11484 3289
rect 11818 3316 13546 3317
rect 11818 3286 12754 3316
rect 11453 3255 11490 3286
rect 9748 3252 11490 3255
rect 1504 3236 1604 3237
rect 2096 2988 2192 3010
rect 1805 2970 1863 2976
rect 1805 2936 1817 2970
rect 1851 2967 1863 2970
rect 2096 2967 2132 2988
rect 1851 2939 2132 2967
rect 1851 2936 1863 2939
rect 1805 2930 1863 2936
rect 2096 2936 2132 2939
rect 2184 2967 2192 2988
rect 2285 2970 2343 2976
rect 2285 2967 2297 2970
rect 2184 2939 2297 2967
rect 2184 2936 2192 2939
rect 2096 2910 2192 2936
rect 2285 2936 2297 2939
rect 2331 2967 2343 2970
rect 2477 2970 2535 2976
rect 2918 2974 2972 3237
rect 3560 3233 5288 3250
rect 2477 2967 2489 2970
rect 2331 2939 2489 2967
rect 2331 2936 2343 2939
rect 2285 2930 2343 2936
rect 2477 2936 2489 2939
rect 2523 2936 2535 2970
rect 2477 2930 2535 2936
rect 2858 2940 2990 2974
rect 2376 2896 2446 2910
rect 2376 2862 2396 2896
rect 2430 2862 2446 2896
rect 2858 2898 2920 2940
rect 2960 2898 2990 2940
rect 3166 2972 3920 2978
rect 3166 2966 3925 2972
rect 3166 2960 3879 2966
rect 3166 2926 3174 2960
rect 3208 2932 3879 2960
rect 3913 2963 3925 2966
rect 4347 2966 4405 2972
rect 4347 2963 4359 2966
rect 3913 2935 4359 2963
rect 3913 2932 3925 2935
rect 3208 2926 3925 2932
rect 4347 2932 4359 2935
rect 4393 2963 4405 2966
rect 4539 2966 4597 2972
rect 4980 2970 5034 3233
rect 5634 3231 7362 3250
rect 5218 2972 5274 3004
rect 5218 2970 5978 2972
rect 4539 2963 4551 2966
rect 4393 2935 4551 2963
rect 4393 2932 4405 2935
rect 4347 2926 4405 2932
rect 4539 2932 4551 2935
rect 4585 2932 4597 2966
rect 4539 2926 4597 2932
rect 4920 2936 5052 2970
rect 3166 2912 3920 2926
rect 2858 2888 2990 2898
rect 4438 2892 4508 2906
rect 2376 2830 2446 2862
rect 4438 2858 4458 2892
rect 4492 2858 4508 2892
rect 4920 2894 4982 2936
rect 5022 2894 5052 2936
rect 5218 2964 5999 2970
rect 5218 2962 5953 2964
rect 5218 2928 5232 2962
rect 5268 2930 5953 2962
rect 5987 2961 5999 2964
rect 6421 2964 6479 2970
rect 6421 2961 6433 2964
rect 5987 2933 6433 2961
rect 5987 2930 5999 2933
rect 5268 2928 5999 2930
rect 5218 2924 5999 2928
rect 6421 2930 6433 2933
rect 6467 2961 6479 2964
rect 6613 2964 6671 2970
rect 7054 2968 7108 3231
rect 7696 3227 9424 3250
rect 9756 3238 11490 3252
rect 11814 3285 12754 3286
rect 12816 3290 13546 3316
rect 13892 3304 15612 3315
rect 13892 3290 14806 3304
rect 12816 3285 13558 3290
rect 11814 3251 11849 3285
rect 11883 3251 11945 3285
rect 11979 3251 12041 3285
rect 12075 3251 12137 3285
rect 12171 3251 12233 3285
rect 12267 3251 12329 3285
rect 12363 3251 12425 3285
rect 12459 3251 12521 3285
rect 12555 3251 12617 3285
rect 12651 3251 12713 3285
rect 12747 3254 12754 3285
rect 12747 3251 12809 3254
rect 12843 3251 12905 3285
rect 12939 3251 13001 3285
rect 13035 3251 13097 3285
rect 13131 3251 13193 3285
rect 13227 3251 13289 3285
rect 13323 3251 13385 3285
rect 13419 3251 13481 3285
rect 13515 3251 13558 3285
rect 11814 3242 13558 3251
rect 13882 3283 14806 3290
rect 14868 3283 15612 3304
rect 15954 3308 17682 3311
rect 15954 3290 16854 3308
rect 13882 3249 13923 3283
rect 13957 3249 14019 3283
rect 14053 3249 14115 3283
rect 14149 3249 14211 3283
rect 14245 3249 14307 3283
rect 14341 3249 14403 3283
rect 14437 3249 14499 3283
rect 14533 3249 14595 3283
rect 14629 3249 14691 3283
rect 14725 3249 14787 3283
rect 14868 3249 14883 3283
rect 14917 3249 14979 3283
rect 15013 3249 15075 3283
rect 15109 3249 15171 3283
rect 15205 3249 15267 3283
rect 15301 3249 15363 3283
rect 15397 3249 15459 3283
rect 15493 3249 15555 3283
rect 15589 3249 15612 3283
rect 13882 3242 14806 3249
rect 14868 3242 15612 3249
rect 15936 3279 16854 3290
rect 16916 3279 17682 3308
rect 15936 3245 15985 3279
rect 16019 3245 16081 3279
rect 16115 3245 16177 3279
rect 16211 3245 16273 3279
rect 16307 3245 16369 3279
rect 16403 3245 16465 3279
rect 16499 3245 16561 3279
rect 16595 3245 16657 3279
rect 16691 3245 16753 3279
rect 16787 3245 16849 3279
rect 16916 3246 16945 3279
rect 16883 3245 16945 3246
rect 16979 3245 17041 3279
rect 17075 3245 17137 3279
rect 17171 3245 17233 3279
rect 17267 3245 17329 3279
rect 17363 3245 17425 3279
rect 17459 3245 17521 3279
rect 17555 3245 17617 3279
rect 17651 3245 17682 3279
rect 15936 3242 17682 3245
rect 11814 3238 13546 3242
rect 6613 2961 6625 2964
rect 6467 2933 6625 2961
rect 6467 2930 6479 2933
rect 6421 2924 6479 2930
rect 6613 2930 6625 2933
rect 6659 2930 6671 2964
rect 6613 2924 6671 2930
rect 6994 2934 7126 2968
rect 5218 2914 5978 2924
rect 5218 2910 5274 2914
rect 4920 2884 5052 2894
rect 6512 2890 6582 2904
rect 2392 2669 2424 2830
rect 4438 2826 4508 2858
rect 6512 2856 6532 2890
rect 6566 2856 6582 2890
rect 6994 2892 7056 2934
rect 7096 2892 7126 2934
rect 7302 2966 8056 2972
rect 7302 2960 8061 2966
rect 7302 2954 8015 2960
rect 7302 2920 7310 2954
rect 7344 2926 8015 2954
rect 8049 2957 8061 2960
rect 8483 2960 8541 2966
rect 8483 2957 8495 2960
rect 8049 2929 8495 2957
rect 8049 2926 8061 2929
rect 7344 2920 8061 2926
rect 8483 2926 8495 2929
rect 8529 2957 8541 2960
rect 8675 2960 8733 2966
rect 9116 2964 9170 3227
rect 9756 3223 11484 3238
rect 8675 2957 8687 2960
rect 8529 2929 8687 2957
rect 8529 2926 8541 2929
rect 8483 2920 8541 2926
rect 8675 2926 8687 2929
rect 8721 2926 8733 2960
rect 8675 2920 8733 2926
rect 9056 2930 9188 2964
rect 9362 2962 10114 2966
rect 7302 2906 8056 2920
rect 6994 2882 7126 2892
rect 8574 2886 8644 2900
rect 1498 2664 3226 2669
rect 4454 2665 4486 2826
rect 6512 2824 6582 2856
rect 8574 2852 8594 2886
rect 8628 2852 8644 2886
rect 9056 2888 9118 2930
rect 9158 2888 9188 2930
rect 9354 2956 10121 2962
rect 9354 2944 10075 2956
rect 9354 2910 9366 2944
rect 9402 2922 10075 2944
rect 10109 2953 10121 2956
rect 10543 2956 10601 2962
rect 10543 2953 10555 2956
rect 10109 2925 10555 2953
rect 10109 2922 10121 2925
rect 9402 2916 10121 2922
rect 10543 2922 10555 2925
rect 10589 2953 10601 2956
rect 10735 2956 10793 2962
rect 11176 2960 11230 3223
rect 11818 3219 13546 3238
rect 10735 2953 10747 2956
rect 10589 2925 10747 2953
rect 10589 2922 10601 2925
rect 10543 2916 10601 2922
rect 10735 2922 10747 2925
rect 10781 2922 10793 2956
rect 10735 2916 10793 2922
rect 11116 2926 11248 2960
rect 9402 2910 10114 2916
rect 9354 2900 10114 2910
rect 9362 2898 10114 2900
rect 9056 2878 9188 2888
rect 10634 2882 10704 2896
rect 1496 2646 3226 2664
rect 1496 2637 2426 2646
rect 2488 2638 3226 2646
rect 3560 2642 5288 2665
rect 6528 2663 6560 2824
rect 8574 2820 8644 2852
rect 10634 2848 10654 2882
rect 10688 2848 10704 2882
rect 11116 2884 11178 2926
rect 11218 2884 11248 2926
rect 11424 2958 12178 2964
rect 11424 2952 12183 2958
rect 11424 2946 12137 2952
rect 11424 2912 11432 2946
rect 11466 2918 12137 2946
rect 12171 2949 12183 2952
rect 12605 2952 12663 2958
rect 12605 2949 12617 2952
rect 12171 2921 12617 2949
rect 12171 2918 12183 2921
rect 11466 2912 12183 2918
rect 12605 2918 12617 2921
rect 12651 2949 12663 2952
rect 12797 2952 12855 2958
rect 13238 2956 13292 3219
rect 13892 3217 15612 3242
rect 13476 2958 13532 2990
rect 13476 2956 14236 2958
rect 12797 2949 12809 2952
rect 12651 2921 12809 2949
rect 12651 2918 12663 2921
rect 12605 2912 12663 2918
rect 12797 2918 12809 2921
rect 12843 2918 12855 2952
rect 12797 2912 12855 2918
rect 13178 2922 13310 2956
rect 11424 2898 12178 2912
rect 11116 2874 11248 2884
rect 12696 2878 12766 2892
rect 5634 2660 7358 2663
rect 5634 2642 6506 2660
rect 3560 2638 5302 2642
rect 2488 2637 3232 2638
rect 1496 2603 1529 2637
rect 1563 2603 1625 2637
rect 1659 2603 1721 2637
rect 1755 2603 1817 2637
rect 1851 2603 1913 2637
rect 1947 2603 2009 2637
rect 2043 2603 2105 2637
rect 2139 2603 2201 2637
rect 2235 2603 2297 2637
rect 2331 2603 2393 2637
rect 2488 2603 2489 2637
rect 2523 2603 2585 2637
rect 2619 2603 2681 2637
rect 2715 2603 2777 2637
rect 2811 2603 2873 2637
rect 2907 2603 2969 2637
rect 3003 2603 3065 2637
rect 3099 2603 3161 2637
rect 3195 2603 3232 2637
rect 1496 2584 2426 2603
rect 2488 2590 3232 2603
rect 3556 2633 4450 2638
rect 4512 2633 5302 2638
rect 3556 2599 3591 2633
rect 3625 2599 3687 2633
rect 3721 2599 3783 2633
rect 3817 2599 3879 2633
rect 3913 2599 3975 2633
rect 4009 2599 4071 2633
rect 4105 2599 4167 2633
rect 4201 2599 4263 2633
rect 4297 2599 4359 2633
rect 4393 2599 4450 2633
rect 4512 2599 4551 2633
rect 4585 2599 4647 2633
rect 4681 2599 4743 2633
rect 4777 2599 4839 2633
rect 4873 2599 4935 2633
rect 4969 2599 5031 2633
rect 5065 2599 5127 2633
rect 5161 2599 5223 2633
rect 5257 2599 5302 2633
rect 3556 2590 4450 2599
rect 2488 2584 3226 2590
rect 1496 2582 3226 2584
rect 1498 2571 3226 2582
rect 3560 2576 4450 2590
rect 4512 2594 5302 2599
rect 5626 2631 6506 2642
rect 6568 2631 7358 2660
rect 8590 2659 8622 2820
rect 10634 2816 10704 2848
rect 12696 2844 12716 2878
rect 12750 2844 12766 2878
rect 13178 2880 13240 2922
rect 13280 2880 13310 2922
rect 13476 2950 14257 2956
rect 13476 2948 14211 2950
rect 13476 2914 13490 2948
rect 13526 2916 14211 2948
rect 14245 2947 14257 2950
rect 14679 2950 14737 2956
rect 14679 2947 14691 2950
rect 14245 2919 14691 2947
rect 14245 2916 14257 2919
rect 13526 2914 14257 2916
rect 13476 2910 14257 2914
rect 14679 2916 14691 2919
rect 14725 2947 14737 2950
rect 14871 2950 14929 2956
rect 15312 2954 15366 3217
rect 15954 3213 17682 3242
rect 14871 2947 14883 2950
rect 14725 2919 14883 2947
rect 14725 2916 14737 2919
rect 14679 2910 14737 2916
rect 14871 2916 14883 2919
rect 14917 2916 14929 2950
rect 14871 2910 14929 2916
rect 15252 2920 15384 2954
rect 13476 2900 14236 2910
rect 13476 2896 13532 2900
rect 13178 2870 13310 2880
rect 14770 2876 14840 2890
rect 5626 2597 5665 2631
rect 5699 2597 5761 2631
rect 5795 2597 5857 2631
rect 5891 2597 5953 2631
rect 5987 2597 6049 2631
rect 6083 2597 6145 2631
rect 6179 2597 6241 2631
rect 6275 2597 6337 2631
rect 6371 2597 6433 2631
rect 6467 2598 6506 2631
rect 6568 2598 6625 2631
rect 6467 2597 6529 2598
rect 6563 2597 6625 2598
rect 6659 2597 6721 2631
rect 6755 2597 6817 2631
rect 6851 2597 6913 2631
rect 6947 2597 7009 2631
rect 7043 2597 7105 2631
rect 7139 2597 7201 2631
rect 7235 2597 7297 2631
rect 7331 2597 7358 2631
rect 7696 2642 9424 2659
rect 10650 2655 10682 2816
rect 12696 2812 12766 2844
rect 14770 2842 14790 2876
rect 14824 2842 14840 2876
rect 15252 2878 15314 2920
rect 15354 2878 15384 2920
rect 15560 2952 16314 2958
rect 15560 2946 16319 2952
rect 15560 2940 16273 2946
rect 15560 2906 15568 2940
rect 15602 2912 16273 2940
rect 16307 2943 16319 2946
rect 16741 2946 16799 2952
rect 16741 2943 16753 2946
rect 16307 2915 16753 2943
rect 16307 2912 16319 2915
rect 15602 2906 16319 2912
rect 16741 2912 16753 2915
rect 16787 2943 16799 2946
rect 16933 2946 16991 2952
rect 17374 2950 17428 3213
rect 16933 2943 16945 2946
rect 16787 2915 16945 2943
rect 16787 2912 16799 2915
rect 16741 2906 16799 2912
rect 16933 2912 16945 2915
rect 16979 2912 16991 2946
rect 16933 2906 16991 2912
rect 17314 2916 17446 2950
rect 15560 2892 16314 2906
rect 15252 2868 15384 2878
rect 16832 2872 16902 2886
rect 7696 2627 8556 2642
rect 8618 2627 9424 2642
rect 7696 2626 7727 2627
rect 5626 2594 7358 2597
rect 4512 2576 5288 2594
rect 3560 2567 5288 2576
rect 5634 2565 7358 2594
rect 7682 2593 7727 2626
rect 7761 2593 7823 2627
rect 7857 2593 7919 2627
rect 7953 2593 8015 2627
rect 8049 2593 8111 2627
rect 8145 2593 8207 2627
rect 8241 2593 8303 2627
rect 8337 2593 8399 2627
rect 8433 2593 8495 2627
rect 8529 2593 8556 2627
rect 8625 2593 8687 2627
rect 8721 2593 8783 2627
rect 8817 2593 8879 2627
rect 8913 2593 8975 2627
rect 9009 2593 9071 2627
rect 9105 2593 9167 2627
rect 9201 2593 9263 2627
rect 9297 2593 9359 2627
rect 9393 2626 9424 2627
rect 9756 2642 11484 2655
rect 12712 2651 12744 2812
rect 14770 2810 14840 2842
rect 16832 2838 16852 2872
rect 16886 2838 16902 2872
rect 17314 2874 17376 2916
rect 17416 2874 17446 2916
rect 17314 2864 17446 2874
rect 17610 2872 17738 2876
rect 9756 2626 10724 2642
rect 9393 2593 9426 2626
rect 7682 2580 8556 2593
rect 8618 2580 9426 2593
rect 7682 2578 9426 2580
rect 9750 2623 10724 2626
rect 10786 2623 11484 2642
rect 9750 2589 9787 2623
rect 9821 2589 9883 2623
rect 9917 2589 9979 2623
rect 10013 2589 10075 2623
rect 10109 2589 10171 2623
rect 10205 2589 10267 2623
rect 10301 2589 10363 2623
rect 10397 2589 10459 2623
rect 10493 2589 10555 2623
rect 10589 2589 10651 2623
rect 10685 2589 10724 2623
rect 10786 2589 10843 2623
rect 10877 2589 10939 2623
rect 10973 2589 11035 2623
rect 11069 2589 11131 2623
rect 11165 2589 11227 2623
rect 11261 2589 11323 2623
rect 11357 2589 11419 2623
rect 11453 2622 11484 2623
rect 11818 2632 13546 2651
rect 14786 2649 14818 2810
rect 16832 2806 16902 2838
rect 17610 2862 17940 2872
rect 17610 2846 17812 2862
rect 17610 2808 17616 2846
rect 17658 2808 17812 2846
rect 11818 2622 12748 2632
rect 11453 2589 11490 2622
rect 9750 2580 10724 2589
rect 10786 2580 11490 2589
rect 9750 2578 11490 2580
rect 7696 2561 9424 2578
rect 9756 2574 11490 2578
rect 11814 2619 12748 2622
rect 12810 2622 13546 2632
rect 13892 2636 15620 2649
rect 16848 2645 16880 2806
rect 17610 2774 17812 2808
rect 17902 2774 17940 2862
rect 17610 2758 17940 2774
rect 13892 2622 14848 2636
rect 12810 2619 13556 2622
rect 11814 2585 11849 2619
rect 11883 2585 11945 2619
rect 11979 2585 12041 2619
rect 12075 2585 12137 2619
rect 12171 2585 12233 2619
rect 12267 2585 12329 2619
rect 12363 2585 12425 2619
rect 12459 2585 12521 2619
rect 12555 2585 12617 2619
rect 12651 2585 12713 2619
rect 12747 2585 12748 2619
rect 12843 2585 12905 2619
rect 12939 2585 13001 2619
rect 13035 2585 13097 2619
rect 13131 2585 13193 2619
rect 13227 2585 13289 2619
rect 13323 2585 13385 2619
rect 13419 2585 13481 2619
rect 13515 2585 13556 2619
rect 11814 2574 12748 2585
rect 9756 2557 11484 2574
rect 11818 2570 12748 2574
rect 12810 2574 13556 2585
rect 13880 2617 14848 2622
rect 14910 2626 15620 2636
rect 15954 2630 17682 2645
rect 15954 2626 16896 2630
rect 14910 2617 15624 2626
rect 13880 2583 13923 2617
rect 13957 2583 14019 2617
rect 14053 2583 14115 2617
rect 14149 2583 14211 2617
rect 14245 2583 14307 2617
rect 14341 2583 14403 2617
rect 14437 2583 14499 2617
rect 14533 2583 14595 2617
rect 14629 2583 14691 2617
rect 14725 2583 14787 2617
rect 14821 2583 14848 2617
rect 14917 2583 14979 2617
rect 15013 2583 15075 2617
rect 15109 2583 15171 2617
rect 15205 2583 15267 2617
rect 15301 2583 15363 2617
rect 15397 2583 15459 2617
rect 15493 2583 15555 2617
rect 15589 2583 15624 2617
rect 13880 2574 14848 2583
rect 14910 2578 15624 2583
rect 15948 2613 16896 2626
rect 16958 2613 17682 2630
rect 15948 2579 15985 2613
rect 16019 2579 16081 2613
rect 16115 2579 16177 2613
rect 16211 2579 16273 2613
rect 16307 2579 16369 2613
rect 16403 2579 16465 2613
rect 16499 2579 16561 2613
rect 16595 2579 16657 2613
rect 16691 2579 16753 2613
rect 16787 2579 16849 2613
rect 16883 2579 16896 2613
rect 16979 2579 17041 2613
rect 17075 2579 17137 2613
rect 17171 2579 17233 2613
rect 17267 2579 17329 2613
rect 17363 2579 17425 2613
rect 17459 2579 17521 2613
rect 17555 2579 17617 2613
rect 17651 2579 17682 2613
rect 15948 2578 16896 2579
rect 14910 2574 15620 2578
rect 12810 2570 13546 2574
rect 11818 2553 13546 2570
rect 13892 2551 15620 2574
rect 15954 2568 16896 2578
rect 16958 2568 17682 2579
rect 15954 2547 17682 2568
rect 30392 174 30508 5738
rect 30390 144 30514 174
rect 30390 68 30408 144
rect 30482 68 30514 144
rect 30390 34 30514 68
<< via1 >>
rect 27662 44952 27722 45014
rect 2198 7234 2256 7296
rect 4396 7200 4454 7262
rect 6422 7228 6480 7290
rect 8496 7234 8554 7296
rect 2202 6552 2260 6614
rect 4396 6506 4454 6568
rect 6436 6536 6494 6598
rect 8520 6550 8578 6612
rect 9498 6562 9550 6614
rect 9196 6282 9254 6344
rect 2202 6028 2260 6090
rect 4404 6054 4462 6116
rect 6460 6030 6518 6092
rect 8526 6018 8584 6080
rect 18232 6161 18284 6172
rect 16928 6090 16988 6152
rect 18232 6127 18243 6161
rect 18243 6127 18277 6161
rect 18277 6127 18284 6161
rect 18232 6120 18284 6127
rect 18854 6106 18906 6158
rect 19468 6096 19526 6152
rect 20182 6096 20240 6152
rect 21114 6082 21172 6138
rect 22168 6078 22222 6136
rect 23444 6094 23500 6148
rect 25196 6084 25248 6136
rect 27032 6113 27086 6144
rect 27032 6092 27057 6113
rect 27057 6092 27086 6113
rect 28838 6095 28892 6126
rect 28838 6074 28863 6095
rect 28863 6074 28892 6095
rect 17302 5700 17354 5752
rect 17416 5696 17468 5748
rect 18236 5617 18290 5630
rect 18236 5583 18243 5617
rect 18243 5583 18277 5617
rect 18277 5583 18290 5617
rect 18236 5570 18290 5583
rect 18858 5556 18912 5616
rect 19484 5550 19542 5604
rect 20180 5532 20242 5588
rect 21092 5538 21154 5594
rect 22200 5524 22252 5576
rect 23466 5526 23522 5582
rect 25160 5534 25212 5586
rect 27048 5535 27057 5564
rect 27057 5535 27091 5564
rect 27091 5535 27104 5564
rect 27048 5508 27104 5535
rect 28854 5517 28863 5546
rect 28863 5517 28897 5546
rect 28897 5517 28910 5546
rect 28854 5490 28910 5517
rect 2302 5366 2360 5428
rect 4336 5378 4394 5440
rect 17208 5418 17268 5480
rect 6390 5354 6448 5416
rect 8504 5346 8562 5408
rect 904 4420 958 4486
rect 8192 4138 8244 4142
rect 8192 4096 8220 4138
rect 8220 4096 8244 4138
rect 8192 4090 8244 4096
rect 8312 4146 8364 4196
rect 8312 4144 8320 4146
rect 8320 4144 8354 4146
rect 8354 4144 8364 4146
rect 344 3740 438 3830
rect 2482 3303 2544 3332
rect 2482 3270 2489 3303
rect 2489 3270 2523 3303
rect 2523 3270 2544 3303
rect 4532 3299 4594 3324
rect 4532 3265 4551 3299
rect 4551 3265 4585 3299
rect 4585 3265 4594 3299
rect 4532 3262 4594 3265
rect 6482 3297 6544 3326
rect 6482 3264 6529 3297
rect 6529 3264 6544 3297
rect 8590 3293 8652 3318
rect 8590 3259 8591 3293
rect 8591 3259 8625 3293
rect 8625 3259 8652 3293
rect 8590 3256 8652 3259
rect 10698 3289 10760 3320
rect 10698 3258 10747 3289
rect 10747 3258 10760 3289
rect 2132 2936 2184 2988
rect 12754 3285 12816 3316
rect 12754 3254 12809 3285
rect 12809 3254 12816 3285
rect 14806 3283 14868 3304
rect 14806 3249 14821 3283
rect 14821 3249 14868 3283
rect 14806 3242 14868 3249
rect 16854 3279 16916 3308
rect 16854 3246 16883 3279
rect 16883 3246 16916 3279
rect 2426 2637 2488 2646
rect 2426 2603 2427 2637
rect 2427 2603 2488 2637
rect 2426 2584 2488 2603
rect 4450 2633 4512 2638
rect 4450 2599 4455 2633
rect 4455 2599 4489 2633
rect 4489 2599 4512 2633
rect 4450 2576 4512 2599
rect 6506 2631 6568 2660
rect 6506 2598 6529 2631
rect 6529 2598 6563 2631
rect 6563 2598 6568 2631
rect 8556 2627 8618 2642
rect 8556 2593 8591 2627
rect 8591 2593 8618 2627
rect 8556 2580 8618 2593
rect 10724 2623 10786 2642
rect 10724 2589 10747 2623
rect 10747 2589 10781 2623
rect 10781 2589 10786 2623
rect 10724 2580 10786 2589
rect 12748 2619 12810 2632
rect 17812 2774 17902 2862
rect 12748 2585 12809 2619
rect 12809 2585 12810 2619
rect 12748 2570 12810 2585
rect 14848 2617 14910 2636
rect 14848 2583 14883 2617
rect 14883 2583 14910 2617
rect 14848 2574 14910 2583
rect 16896 2613 16958 2630
rect 16896 2579 16945 2613
rect 16945 2579 16958 2613
rect 16896 2568 16958 2579
rect 30408 68 30482 144
<< metal2 >>
rect 27624 45014 27752 45042
rect 27624 44952 27662 45014
rect 27722 44952 27752 45014
rect 27624 44946 27752 44952
rect 2124 7296 2318 7298
rect 8426 7296 8620 7304
rect 2124 7234 2198 7296
rect 2256 7234 2318 7296
rect 6352 7290 6546 7296
rect 2124 7206 2318 7234
rect 4326 7262 4520 7266
rect 4326 7200 4396 7262
rect 4454 7200 4520 7262
rect 6352 7228 6422 7290
rect 6480 7228 6546 7290
rect 6352 7204 6546 7228
rect 8426 7234 8496 7296
rect 8554 7234 8620 7296
rect 8426 7212 8620 7234
rect 4326 7174 4520 7200
rect 2150 6614 2322 6626
rect 2150 6552 2202 6614
rect 2260 6552 2322 6614
rect 6398 6598 6564 6626
rect 2150 6538 2322 6552
rect 4344 6568 4510 6598
rect 4344 6506 4396 6568
rect 4454 6506 4510 6568
rect 6398 6536 6436 6598
rect 6494 6536 6564 6598
rect 6398 6526 6564 6536
rect 8474 6612 8640 6630
rect 8474 6550 8520 6612
rect 8578 6550 8640 6612
rect 8474 6530 8640 6550
rect 9468 6614 17404 6668
rect 9468 6562 9498 6614
rect 9550 6562 17404 6614
rect 9468 6506 17404 6562
rect 4344 6498 4510 6506
rect 9182 6344 9266 6384
rect 9182 6282 9196 6344
rect 9254 6282 9266 6344
rect 9182 6232 9266 6282
rect 16914 6152 17002 6166
rect 4346 6116 4512 6140
rect 2152 6090 2318 6116
rect 2152 6028 2202 6090
rect 2260 6028 2318 6090
rect 4346 6054 4404 6116
rect 4462 6054 4512 6116
rect 4346 6040 4512 6054
rect 6398 6092 6564 6122
rect 2152 6016 2318 6028
rect 6398 6030 6460 6092
rect 6518 6030 6564 6092
rect 6398 6022 6564 6030
rect 8474 6080 8640 6100
rect 8474 6018 8526 6080
rect 8584 6018 8640 6080
rect 16914 6090 16928 6152
rect 16988 6090 17002 6152
rect 16914 6060 17002 6090
rect 8474 6000 8640 6018
rect 17292 5860 17400 6506
rect 18158 6176 18364 6182
rect 18158 6120 18232 6176
rect 18290 6120 18364 6176
rect 18158 6096 18364 6120
rect 18780 6162 18986 6168
rect 18780 6106 18854 6162
rect 18912 6106 18986 6162
rect 18780 6082 18986 6106
rect 19392 6152 19598 6172
rect 19392 6096 19468 6152
rect 19526 6096 19598 6152
rect 19392 6086 19598 6096
rect 20108 6152 20314 6168
rect 20108 6096 20182 6152
rect 20240 6096 20314 6152
rect 23318 6150 23610 6154
rect 20108 6082 20314 6096
rect 21048 6138 21254 6150
rect 21048 6082 21114 6138
rect 21172 6082 21254 6138
rect 21048 6064 21254 6082
rect 22044 6136 22336 6142
rect 22044 6078 22168 6136
rect 22226 6078 22336 6136
rect 23318 6094 23444 6150
rect 23500 6094 23610 6150
rect 27022 6148 27100 6158
rect 27022 6146 27032 6148
rect 23318 6086 23610 6094
rect 25068 6140 25360 6142
rect 22044 6074 22336 6078
rect 25068 6084 25196 6140
rect 25252 6084 25360 6140
rect 25068 6074 25360 6084
rect 26896 6092 27032 6146
rect 27088 6146 27100 6148
rect 27088 6092 27188 6146
rect 28828 6130 28906 6140
rect 28828 6128 28838 6130
rect 26896 6078 27188 6092
rect 28702 6074 28838 6128
rect 28894 6128 28906 6130
rect 28894 6074 28994 6128
rect 28702 6060 28994 6074
rect 17292 5752 17374 5860
rect 17292 5700 17302 5752
rect 17354 5700 17374 5752
rect 17292 5686 17374 5700
rect 17406 5748 17510 5760
rect 17406 5696 17416 5748
rect 17468 5696 17510 5748
rect 17180 5480 17330 5496
rect 2248 5428 2442 5444
rect 2248 5366 2302 5428
rect 2360 5366 2442 5428
rect 4266 5440 4460 5462
rect 4266 5378 4336 5440
rect 4394 5378 4460 5440
rect 4266 5370 4460 5378
rect 6326 5416 6520 5428
rect 2248 5352 2442 5366
rect 6326 5354 6390 5416
rect 6448 5354 6520 5416
rect 17180 5418 17208 5480
rect 17268 5418 17330 5480
rect 6326 5336 6520 5354
rect 8446 5408 8640 5414
rect 8446 5346 8504 5408
rect 8562 5346 8640 5408
rect 17180 5396 17330 5418
rect 8446 5322 8640 5346
rect 890 4486 972 4516
rect 890 4420 904 4486
rect 960 4420 972 4486
rect 890 4386 972 4420
rect 17406 4262 17510 5696
rect 18124 5630 18372 5644
rect 18124 5570 18236 5630
rect 18292 5570 18372 5630
rect 18124 5548 18372 5570
rect 18746 5616 18994 5630
rect 18746 5556 18858 5616
rect 18914 5556 18994 5616
rect 18746 5534 18994 5556
rect 19378 5606 19626 5628
rect 19378 5550 19484 5606
rect 19542 5550 19626 5606
rect 19378 5532 19626 5550
rect 20070 5588 20318 5628
rect 20070 5532 20180 5588
rect 20242 5532 20318 5588
rect 21014 5594 21262 5600
rect 21014 5538 21092 5594
rect 21154 5538 21262 5594
rect 25044 5592 25334 5606
rect 21014 5504 21262 5538
rect 22082 5580 22374 5592
rect 22082 5524 22200 5580
rect 22256 5524 22374 5580
rect 23362 5582 23654 5588
rect 23362 5526 23466 5582
rect 23522 5526 23654 5582
rect 23362 5520 23654 5526
rect 25044 5534 25160 5592
rect 25216 5572 25334 5592
rect 25216 5534 25336 5572
rect 25044 5504 25336 5534
rect 26910 5564 27202 5572
rect 26910 5508 27048 5564
rect 27104 5508 27202 5564
rect 26910 5504 27202 5508
rect 28716 5546 29008 5554
rect 28716 5490 28854 5546
rect 28910 5490 29008 5546
rect 28716 5486 29008 5490
rect 8297 4196 17922 4262
rect 2126 4142 8254 4174
rect 2126 4090 8192 4142
rect 8244 4090 8254 4142
rect 8297 4144 8312 4196
rect 8364 4144 17922 4196
rect 8297 4128 17922 4144
rect 2126 4070 8254 4090
rect 2126 4044 2244 4070
rect 294 3830 484 3880
rect 294 3740 344 3830
rect 438 3740 484 3830
rect 294 3684 484 3740
rect 2128 2994 2188 4044
rect 2390 3332 2648 3336
rect 2390 3270 2482 3332
rect 2544 3270 2648 3332
rect 2390 3262 2648 3270
rect 4444 3324 4702 3328
rect 4444 3262 4532 3324
rect 4594 3262 4702 3324
rect 6392 3326 6650 3338
rect 6392 3264 6482 3326
rect 6544 3264 6650 3326
rect 10610 3320 10868 3328
rect 8498 3318 8756 3320
rect 4444 3254 4702 3262
rect 8498 3256 8590 3318
rect 8652 3256 8756 3318
rect 8498 3246 8756 3256
rect 10610 3258 10698 3320
rect 10760 3258 10868 3320
rect 10610 3254 10868 3258
rect 12652 3254 12754 3316
rect 12816 3254 12910 3316
rect 12652 3242 12910 3254
rect 14702 3304 14960 3310
rect 14702 3242 14806 3304
rect 14868 3242 14960 3304
rect 14702 3236 14960 3242
rect 16770 3308 17028 3314
rect 16770 3246 16854 3308
rect 16916 3246 17028 3308
rect 16770 3240 17028 3246
rect 2104 2988 2194 2994
rect 2104 2936 2132 2988
rect 2184 2936 2194 2988
rect 2104 2922 2194 2936
rect 17788 2862 17922 4128
rect 17788 2774 17812 2862
rect 17902 2774 17922 2862
rect 6416 2660 6674 2662
rect 2348 2646 2606 2650
rect 2348 2584 2426 2646
rect 2488 2584 2606 2646
rect 2348 2576 2606 2584
rect 4364 2638 4622 2642
rect 4364 2576 4450 2638
rect 4512 2576 4622 2638
rect 6416 2598 6506 2660
rect 6568 2598 6674 2660
rect 6416 2588 6674 2598
rect 8464 2642 8722 2646
rect 4364 2568 4622 2576
rect 8464 2580 8556 2642
rect 8618 2580 8722 2642
rect 8464 2572 8722 2580
rect 10636 2642 10894 2646
rect 10636 2580 10724 2642
rect 10786 2580 10894 2642
rect 10636 2572 10894 2580
rect 12648 2632 12906 2638
rect 12648 2570 12748 2632
rect 12810 2570 12906 2632
rect 12648 2564 12906 2570
rect 14736 2636 14994 2642
rect 14736 2574 14848 2636
rect 14910 2574 14994 2636
rect 14736 2568 14994 2574
rect 16792 2630 17050 2640
rect 16792 2568 16896 2630
rect 16958 2568 17050 2630
rect 16792 2566 17050 2568
rect 30390 144 30514 174
rect 30390 68 30408 144
rect 30482 68 30514 144
rect 30390 34 30514 68
<< via2 >>
rect 27662 44952 27722 45014
rect 2198 7234 2256 7296
rect 4396 7200 4454 7262
rect 6422 7228 6480 7290
rect 8496 7234 8554 7296
rect 2202 6552 2260 6614
rect 4396 6506 4454 6568
rect 6436 6536 6494 6598
rect 8520 6550 8578 6612
rect 9196 6282 9254 6344
rect 2202 6028 2260 6090
rect 4404 6054 4462 6116
rect 6460 6030 6518 6092
rect 8526 6018 8584 6080
rect 16928 6090 16988 6152
rect 18232 6172 18290 6176
rect 18232 6120 18284 6172
rect 18284 6120 18290 6172
rect 18854 6158 18912 6162
rect 18854 6106 18906 6158
rect 18906 6106 18912 6158
rect 19468 6096 19526 6152
rect 20182 6096 20240 6152
rect 21114 6082 21172 6138
rect 22168 6078 22222 6136
rect 22222 6078 22226 6136
rect 23444 6148 23500 6150
rect 23444 6094 23500 6148
rect 25196 6136 25252 6140
rect 25196 6084 25248 6136
rect 25248 6084 25252 6136
rect 27032 6144 27088 6148
rect 27032 6092 27086 6144
rect 27086 6092 27088 6144
rect 28838 6126 28894 6130
rect 28838 6074 28892 6126
rect 28892 6074 28894 6126
rect 2302 5366 2360 5428
rect 4336 5378 4394 5440
rect 6390 5354 6448 5416
rect 17208 5418 17268 5480
rect 8504 5346 8562 5408
rect 904 4420 958 4486
rect 958 4420 960 4486
rect 18236 5570 18290 5630
rect 18290 5570 18292 5630
rect 18858 5556 18912 5616
rect 18912 5556 18914 5616
rect 19484 5604 19542 5606
rect 19484 5550 19542 5604
rect 20180 5532 20242 5588
rect 21092 5538 21154 5594
rect 22200 5576 22256 5580
rect 22200 5524 22252 5576
rect 22252 5524 22256 5576
rect 23466 5526 23522 5582
rect 25160 5586 25216 5592
rect 25160 5534 25212 5586
rect 25212 5534 25216 5586
rect 27048 5508 27104 5564
rect 28854 5490 28910 5546
rect 344 3740 438 3830
rect 2482 3270 2544 3332
rect 4532 3262 4594 3324
rect 6482 3264 6544 3326
rect 8590 3256 8652 3318
rect 10698 3258 10760 3320
rect 12754 3254 12816 3316
rect 14806 3242 14868 3304
rect 16854 3246 16916 3308
rect 2426 2584 2488 2646
rect 4450 2576 4512 2638
rect 6506 2598 6568 2660
rect 8556 2580 8618 2642
rect 10724 2580 10786 2642
rect 12748 2570 12810 2632
rect 14848 2574 14910 2636
rect 16896 2568 16958 2630
rect 30408 68 30482 144
<< metal3 >>
rect 27624 45022 27752 45042
rect 27624 45014 27668 45022
rect 27624 44952 27662 45014
rect 27732 44958 27752 45022
rect 27722 44952 27752 44958
rect 27624 44946 27752 44952
rect 390 7512 9404 7542
rect 390 7386 422 7512
rect 548 7386 9404 7512
rect 390 7340 9404 7386
rect 2123 7296 2325 7340
rect 2123 7234 2198 7296
rect 2256 7234 2325 7296
rect 2123 7215 2325 7234
rect 4323 7262 4525 7340
rect 4323 7200 4396 7262
rect 4454 7200 4525 7262
rect 6345 7290 6547 7340
rect 6345 7228 6422 7290
rect 6480 7228 6547 7290
rect 6345 7209 6547 7228
rect 8429 7296 8631 7340
rect 8429 7234 8496 7296
rect 8554 7234 8631 7296
rect 8429 7209 8631 7234
rect 4323 7179 4525 7200
rect 2150 6614 2326 6638
rect 2150 6552 2202 6614
rect 2260 6552 2326 6614
rect 6394 6598 6570 6626
rect 2150 6396 2326 6552
rect 4342 6568 4518 6590
rect 4342 6506 4396 6568
rect 4454 6506 4518 6568
rect 4342 6396 4518 6506
rect 6394 6536 6436 6598
rect 6494 6536 6570 6598
rect 6394 6396 6570 6536
rect 8470 6612 8646 6634
rect 8470 6550 8520 6612
rect 8578 6550 8646 6612
rect 16797 6608 16999 6617
rect 8470 6396 8646 6550
rect 16779 6408 29620 6608
rect 16779 6406 29619 6408
rect 1020 6350 9290 6396
rect 1020 6260 1068 6350
rect 1160 6344 9290 6350
rect 1160 6282 9196 6344
rect 9254 6282 9290 6344
rect 1160 6260 9290 6282
rect 1020 6220 9290 6260
rect 2150 6090 2326 6220
rect 2150 6028 2202 6090
rect 2260 6028 2326 6090
rect 4342 6116 4518 6220
rect 4342 6054 4404 6116
rect 4462 6054 4518 6116
rect 4342 6036 4518 6054
rect 6394 6092 6570 6220
rect 2150 6016 2326 6028
rect 6394 6030 6460 6092
rect 6518 6030 6570 6092
rect 6394 6012 6570 6030
rect 8470 6080 8646 6220
rect 8470 6018 8526 6080
rect 8584 6018 8646 6080
rect 8470 5998 8646 6018
rect 16797 6152 16999 6406
rect 16797 6090 16928 6152
rect 16988 6090 16999 6152
rect 18169 6176 18371 6406
rect 18169 6120 18232 6176
rect 18290 6120 18371 6176
rect 18169 6099 18371 6120
rect 18791 6162 18993 6406
rect 18791 6106 18854 6162
rect 18912 6106 18993 6162
rect 2243 5428 2445 5449
rect 2243 5366 2302 5428
rect 2360 5366 2445 5428
rect 2243 5154 2445 5366
rect 4265 5440 4467 5459
rect 4265 5378 4336 5440
rect 4394 5378 4467 5440
rect 4265 5154 4467 5378
rect 6325 5416 6527 5425
rect 6325 5354 6390 5416
rect 6448 5354 6527 5416
rect 6325 5154 6527 5354
rect 8447 5408 8649 5437
rect 8447 5346 8504 5408
rect 8562 5346 8649 5408
rect 8447 5154 8649 5346
rect 378 5120 9392 5154
rect 378 4994 422 5120
rect 548 4994 9392 5120
rect 378 4952 9392 4994
rect 890 4486 972 4516
rect 890 4420 904 4486
rect 968 4420 972 4486
rect 890 4386 972 4420
rect 294 3830 484 3880
rect 294 3740 344 3830
rect 438 3740 484 3830
rect 294 3684 484 3740
rect 16797 3608 16999 6090
rect 18791 6085 18993 6106
rect 19381 6152 19583 6406
rect 19381 6096 19468 6152
rect 19526 6096 19583 6152
rect 19381 6077 19583 6096
rect 20115 6357 29619 6406
rect 20115 6152 20317 6357
rect 20115 6096 20182 6152
rect 20240 6096 20317 6152
rect 20115 6069 20317 6096
rect 21041 6138 21243 6357
rect 21041 6082 21114 6138
rect 21172 6082 21243 6138
rect 21041 6055 21243 6082
rect 22104 6136 22304 6357
rect 22104 6078 22168 6136
rect 22226 6078 22304 6136
rect 22104 6034 22304 6078
rect 23380 6150 23580 6357
rect 25114 6158 25314 6357
rect 26946 6166 27146 6357
rect 23380 6094 23444 6150
rect 23500 6094 23580 6150
rect 23380 6074 23580 6094
rect 25066 6140 25362 6158
rect 25066 6084 25196 6140
rect 25252 6084 25362 6140
rect 25066 6074 25362 6084
rect 26892 6148 27190 6166
rect 28752 6148 28952 6357
rect 26892 6092 27032 6148
rect 27088 6092 27190 6148
rect 26892 6072 27190 6092
rect 28698 6130 28996 6148
rect 28698 6074 28838 6130
rect 28894 6074 28996 6130
rect 26946 6052 27146 6072
rect 28698 6054 28996 6074
rect 28752 6034 28952 6054
rect 18071 5630 18369 5641
rect 18071 5570 18236 5630
rect 18292 5570 18369 5630
rect 17179 5480 17549 5539
rect 17179 5418 17208 5480
rect 17268 5418 17549 5480
rect 17179 5338 17549 5418
rect 18071 5352 18369 5570
rect 18693 5616 18991 5627
rect 18693 5556 18858 5616
rect 18914 5556 18991 5616
rect 18064 5338 18450 5352
rect 18693 5338 18991 5556
rect 19349 5606 19647 5625
rect 19349 5550 19484 5606
rect 19542 5550 19647 5606
rect 19349 5338 19647 5550
rect 20043 5588 20341 5613
rect 20043 5532 20180 5588
rect 20242 5532 20341 5588
rect 20043 5338 20341 5532
rect 20983 5594 21281 5603
rect 20983 5538 21092 5594
rect 21154 5538 21281 5594
rect 20983 5338 21281 5538
rect 22077 5580 22375 5593
rect 22077 5524 22200 5580
rect 22256 5524 22375 5580
rect 22077 5338 22375 5524
rect 23353 5582 23651 5614
rect 23353 5526 23466 5582
rect 23522 5526 23651 5582
rect 23353 5338 23651 5526
rect 25043 5592 25341 5601
rect 25043 5534 25160 5592
rect 25216 5534 25341 5592
rect 25043 5338 25341 5534
rect 26909 5564 27207 5601
rect 26909 5508 27048 5564
rect 27104 5508 27207 5564
rect 26909 5338 27207 5508
rect 28715 5546 29013 5583
rect 28715 5490 28854 5546
rect 28910 5490 29013 5546
rect 28715 5338 29013 5490
rect 17179 5336 20428 5338
rect 20983 5336 28595 5338
rect 17179 5332 28595 5336
rect 28715 5332 29657 5338
rect 17179 4968 29657 5332
rect 464 3566 17010 3608
rect 464 3500 508 3566
rect 572 3500 17010 3566
rect 464 3450 17010 3500
rect 524 3428 17010 3450
rect 1504 3406 17010 3428
rect 2401 3332 2603 3406
rect 2401 3270 2482 3332
rect 2544 3270 2603 3332
rect 2401 3209 2603 3270
rect 4449 3324 4651 3406
rect 4449 3262 4532 3324
rect 4594 3262 4651 3324
rect 4449 3243 4651 3262
rect 6417 3326 6619 3406
rect 6417 3264 6482 3326
rect 6544 3264 6619 3326
rect 6417 3243 6619 3264
rect 8509 3318 8711 3406
rect 8509 3256 8590 3318
rect 8652 3256 8711 3318
rect 8509 3243 8711 3256
rect 10645 3320 10847 3406
rect 10645 3258 10698 3320
rect 10760 3258 10847 3320
rect 10645 3223 10847 3258
rect 12687 3316 12889 3406
rect 12687 3254 12754 3316
rect 12816 3254 12889 3316
rect 12687 3243 12889 3254
rect 14731 3304 14933 3406
rect 14731 3242 14806 3304
rect 14868 3242 14933 3304
rect 14731 3211 14933 3242
rect 16797 3308 16999 3406
rect 16797 3246 16854 3308
rect 16916 3246 16999 3308
rect 16797 3223 16999 3246
rect 2352 2646 2612 2692
rect 2352 2584 2426 2646
rect 2488 2584 2612 2646
rect 2352 2266 2612 2584
rect 4356 2638 4616 2692
rect 4356 2576 4450 2638
rect 4512 2576 4616 2638
rect 4356 2266 4616 2576
rect 6418 2660 6678 2692
rect 6418 2598 6506 2660
rect 6568 2598 6678 2660
rect 6418 2266 6678 2598
rect 8466 2642 8726 2660
rect 8466 2580 8556 2642
rect 8618 2580 8726 2642
rect 8466 2266 8726 2580
rect 10628 2642 10888 2648
rect 10628 2580 10724 2642
rect 10786 2580 10888 2642
rect 10628 2266 10888 2580
rect 12646 2632 12906 2642
rect 12646 2570 12748 2632
rect 12810 2570 12906 2632
rect 12646 2266 12906 2570
rect 14732 2636 14992 2642
rect 14732 2574 14848 2636
rect 14910 2574 14992 2636
rect 14732 2266 14992 2574
rect 16780 2630 17040 2636
rect 16780 2568 16896 2630
rect 16958 2568 17040 2630
rect 16780 2266 17040 2568
rect 17223 2266 17521 4968
rect 1006 2154 17558 2266
rect 1006 2052 1048 2154
rect 1146 2052 17558 2154
rect 1006 1968 17558 2052
rect 30390 144 30514 174
rect 30390 68 30408 144
rect 30482 68 30514 144
rect 30390 34 30514 68
<< via3 >>
rect 27668 45014 27732 45022
rect 27668 44958 27722 45014
rect 27722 44958 27732 45014
rect 422 7386 548 7512
rect 1068 6260 1160 6350
rect 422 4994 548 5120
rect 904 4420 960 4486
rect 960 4420 968 4486
rect 344 3740 438 3830
rect 508 3500 572 3566
rect 1048 2052 1146 2154
rect 30408 68 30482 144
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 45026 27722 45152
rect 27662 45022 27734 45026
rect 27662 44958 27668 45022
rect 27732 44958 27734 45022
rect 27662 44956 27734 44958
rect 27662 44952 27722 44956
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 7512 600 44152
rect 200 7386 422 7512
rect 548 7386 600 7512
rect 200 5120 600 7386
rect 200 4994 422 5120
rect 548 4994 600 5120
rect 200 3830 600 4994
rect 200 3740 344 3830
rect 438 3740 600 3830
rect 200 3566 600 3740
rect 200 3500 508 3566
rect 572 3500 600 3566
rect 200 1000 600 3500
rect 800 6350 1200 44152
rect 800 6260 1068 6350
rect 1160 6260 1200 6350
rect 800 4486 1200 6260
rect 800 4420 904 4486
rect 968 4420 1200 4486
rect 800 2154 1200 4420
rect 800 2052 1048 2154
rect 1146 2052 1200 2154
rect 800 1000 1200 2052
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 144 30542 200
rect 30362 68 30408 144
rect 30482 68 30542 144
rect 30362 0 30542 68
use inverter  inverter_0
timestamp 1752867815
transform -1 0 9366 0 -1 6069
box -578 -1231 8018 743
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1752700594
transform 1 0 18744 0 1 5586
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1752700594
transform 1 0 18122 0 1 5600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1752700594
transform 1 0 19368 0 1 5584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1752700594
transform 1 0 19976 0 1 5572
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  sky130_fd_sc_hd__inv_6_0 pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1752700594
transform 1 0 20800 0 1 5558
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1752774549
transform 1 0 21782 0 1 5562
box -38 -48 866 592
use sky130_fd_sc_hd__inv_12  sky130_fd_sc_hd__inv_12_0 pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1752774549
transform 1 0 22946 0 1 5562
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1752774389
transform 1 0 24476 0 1 5552
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1752774389
transform 1 0 26292 0 1 5552
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1752774389
transform 1 0 28098 0 1 5534
box -38 -48 1510 592
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_0 pdks/sky130B/libs.ref/sky130_fd_sc_hs/mag
timestamp 1752867815
transform 1 0 1498 0 1 2620
box -38 -49 1766 715
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_1
timestamp 1752867815
transform 1 0 3560 0 1 2616
box -38 -49 1766 715
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_2
timestamp 1752867815
transform 1 0 7696 0 1 2610
box -38 -49 1766 715
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_3
timestamp 1752867815
transform 1 0 5634 0 1 2614
box -38 -49 1766 715
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_4
timestamp 1752867815
transform 1 0 13892 0 1 2600
box -38 -49 1766 715
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_5
timestamp 1752867815
transform 1 0 15954 0 1 2596
box -38 -49 1766 715
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_6
timestamp 1752867815
transform 1 0 11818 0 1 2602
box -38 -49 1766 715
use sky130_fd_sc_hs__fa_1  sky130_fd_sc_hs__fa_1_7
timestamp 1752867815
transform 1 0 9756 0 1 2606
box -38 -49 1766 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_0 pdks/sky130B/libs.ref/sky130_fd_sc_hs/mag
timestamp 1752773148
transform -1 0 8386 0 -1 4452
box -38 -49 326 715
use sky130_fd_sc_hs__mux2_1  sky130_fd_sc_hs__mux2_1_0 pdks/sky130B/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 16918 0 1 5448
box -38 -49 902 715
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel comment s 3560 2616 3560 2616 4 fa_1
flabel pwell s 3560 2616 5288 2665 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 3560 3233 5288 3282 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 3560 3233 5288 3282 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 3560 2616 5288 2665 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 4455 2858 4489 2892 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 4935 2932 4969 2966 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 3591 2710 3625 2744 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 3591 2784 3625 2818 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 1498 2620 1498 2620 4 fa_1
flabel pwell s 1498 2620 3226 2669 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 1498 3237 3226 3286 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 2297 2936 2331 2970 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel metal1 s 1498 3237 3226 3286 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 1498 2620 3226 2669 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2393 2862 2427 2896 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2873 2936 2907 2970 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1529 2714 1563 2748 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1529 2788 1563 2822 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 5665 2782 5699 2816 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 5665 2708 5699 2742 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 7009 2930 7043 2964 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 6529 2856 6563 2890 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 5634 2614 7362 2663 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 5634 3231 7362 3280 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel nwell s 5634 3231 7362 3280 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 5634 2614 7362 2663 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 5634 2614 5634 2614 4 fa_1
flabel locali s 7727 2778 7761 2812 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 7727 2704 7761 2738 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 9071 2926 9105 2960 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 8591 2852 8625 2886 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 7696 2610 9424 2659 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 7696 3227 9424 3276 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel nwell s 7696 3227 9424 3276 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 7696 2610 9424 2659 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 7696 2610 7696 2610 4 fa_1
rlabel comment s 13892 2600 13892 2600 4 fa_1
flabel pwell s 13892 2600 15620 2649 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 13892 3217 15620 3266 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 13892 3217 15620 3266 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 13892 2600 15620 2649 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 14787 2842 14821 2876 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 15267 2916 15301 2950 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 13923 2694 13957 2728 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 13923 2768 13957 2802 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 15954 2596 15954 2596 4 fa_1
flabel pwell s 15954 2596 17682 2645 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 15954 3213 17682 3262 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 15954 3213 17682 3262 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 15954 2596 17682 2645 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 16849 2838 16883 2872 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 17329 2912 17363 2946 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 17617 2690 17651 2724 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2764 17651 2798 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2838 17651 2872 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2912 17651 2946 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2986 17651 3020 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 3060 17651 3094 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 3134 17651 3168 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 15985 2690 16019 2724 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 15985 2764 16019 2798 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 11818 2602 11818 2602 4 fa_1
flabel pwell s 11818 2602 13546 2651 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 11818 3219 13546 3268 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 11818 3219 13546 3268 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 11818 2602 13546 2651 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 12713 2844 12747 2878 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 13193 2918 13227 2952 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 11849 2696 11883 2730 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 11849 2770 11883 2804 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 9756 2606 9756 2606 4 fa_1
flabel pwell s 9756 2606 11484 2655 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 9756 3223 11484 3272 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 9756 3223 11484 3272 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 9756 2606 11484 2655 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 10651 2848 10685 2882 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 11131 2922 11165 2956 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 9787 2700 9821 2734 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 9787 2774 9821 2808 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
