magic
tech sky130B
magscale 1 2
timestamp 1752698750
<< nwell >>
rect 8060 3748 8424 4120
rect 1460 2952 3264 3324
rect 1798 2931 2994 2952
rect 3522 2948 5326 3320
rect 3860 2927 5056 2948
rect 5596 2946 7400 3318
rect 5934 2925 7130 2946
rect 7658 2942 9462 3314
rect 7996 2921 9192 2942
rect 9718 2938 11522 3310
rect 10056 2917 11252 2938
rect 11780 2934 13584 3306
rect 12118 2913 13314 2934
rect 13854 2932 15658 3304
rect 14192 2911 15388 2932
rect 15916 2928 17720 3300
rect 16254 2907 17450 2928
rect 22506 2847 22858 3168
rect 23130 2845 23482 3166
rect 23738 2833 24274 3154
rect 24562 2819 25282 3140
<< pwell >>
rect 8098 4403 8386 4452
rect 8100 4204 8382 4403
rect 1499 2849 1688 2868
rect 3036 2849 3225 2868
rect 1499 2669 3225 2849
rect 3561 2845 3750 2864
rect 5098 2845 5287 2864
rect 1498 2620 3226 2669
rect 3561 2665 5287 2845
rect 5635 2843 5824 2862
rect 7172 2843 7361 2862
rect 3560 2616 5288 2665
rect 5635 2663 7361 2843
rect 7697 2839 7886 2858
rect 9234 2839 9423 2858
rect 5634 2614 7362 2663
rect 7697 2659 9423 2839
rect 9757 2835 9946 2854
rect 11294 2835 11483 2854
rect 7696 2610 9424 2659
rect 9757 2655 11483 2835
rect 11819 2831 12008 2850
rect 13356 2831 13545 2850
rect 9756 2606 11484 2655
rect 11819 2651 13545 2831
rect 13893 2829 14082 2848
rect 15430 2829 15619 2848
rect 11818 2602 13546 2651
rect 13893 2649 15619 2829
rect 15955 2825 16144 2844
rect 17492 2825 17681 2844
rect 13892 2600 15620 2649
rect 15955 2645 17681 2825
rect 15954 2596 17682 2645
rect 22586 2607 22772 2789
rect 22586 2603 22607 2607
rect 23171 2605 23441 2787
rect 22573 2569 22607 2603
rect 23197 2567 23231 2605
rect 23787 2593 24225 2775
rect 23805 2555 23839 2593
rect 24611 2579 25243 2761
rect 24629 2541 24663 2579
<< scnmos >>
rect 22664 2633 22694 2763
rect 23249 2631 23279 2761
rect 23333 2631 23363 2761
rect 23865 2619 23895 2749
rect 23949 2619 23979 2749
rect 24033 2619 24063 2749
rect 24117 2619 24147 2749
rect 24713 2605 24743 2735
rect 24797 2605 24827 2735
rect 24881 2605 24911 2735
rect 24965 2605 24995 2735
rect 25049 2605 25079 2735
rect 25133 2605 25163 2735
<< scpmos >>
rect 8182 3860 8212 4084
rect 8272 3860 8302 4084
rect 1582 2988 1612 3212
rect 1685 2988 1715 3188
rect 1786 3009 1816 3209
rect 1887 2967 1917 3167
rect 1977 2967 2007 3167
rect 2074 2967 2104 3167
rect 2191 2967 2221 3167
rect 2292 2967 2322 3167
rect 2384 2967 2414 3167
rect 2485 2967 2515 3167
rect 2575 2967 2605 3167
rect 2694 2967 2724 3167
rect 2861 2982 2891 3182
rect 3112 2988 3142 3212
rect 3644 2984 3674 3208
rect 3747 2984 3777 3184
rect 3848 3005 3878 3205
rect 3949 2963 3979 3163
rect 4039 2963 4069 3163
rect 4136 2963 4166 3163
rect 4253 2963 4283 3163
rect 4354 2963 4384 3163
rect 4446 2963 4476 3163
rect 4547 2963 4577 3163
rect 4637 2963 4667 3163
rect 4756 2963 4786 3163
rect 4923 2978 4953 3178
rect 5174 2984 5204 3208
rect 5718 2982 5748 3206
rect 5821 2982 5851 3182
rect 5922 3003 5952 3203
rect 6023 2961 6053 3161
rect 6113 2961 6143 3161
rect 6210 2961 6240 3161
rect 6327 2961 6357 3161
rect 6428 2961 6458 3161
rect 6520 2961 6550 3161
rect 6621 2961 6651 3161
rect 6711 2961 6741 3161
rect 6830 2961 6860 3161
rect 6997 2976 7027 3176
rect 7248 2982 7278 3206
rect 7780 2978 7810 3202
rect 7883 2978 7913 3178
rect 7984 2999 8014 3199
rect 8085 2957 8115 3157
rect 8175 2957 8205 3157
rect 8272 2957 8302 3157
rect 8389 2957 8419 3157
rect 8490 2957 8520 3157
rect 8582 2957 8612 3157
rect 8683 2957 8713 3157
rect 8773 2957 8803 3157
rect 8892 2957 8922 3157
rect 9059 2972 9089 3172
rect 9310 2978 9340 3202
rect 9840 2974 9870 3198
rect 9943 2974 9973 3174
rect 10044 2995 10074 3195
rect 10145 2953 10175 3153
rect 10235 2953 10265 3153
rect 10332 2953 10362 3153
rect 10449 2953 10479 3153
rect 10550 2953 10580 3153
rect 10642 2953 10672 3153
rect 10743 2953 10773 3153
rect 10833 2953 10863 3153
rect 10952 2953 10982 3153
rect 11119 2968 11149 3168
rect 11370 2974 11400 3198
rect 11902 2970 11932 3194
rect 12005 2970 12035 3170
rect 12106 2991 12136 3191
rect 12207 2949 12237 3149
rect 12297 2949 12327 3149
rect 12394 2949 12424 3149
rect 12511 2949 12541 3149
rect 12612 2949 12642 3149
rect 12704 2949 12734 3149
rect 12805 2949 12835 3149
rect 12895 2949 12925 3149
rect 13014 2949 13044 3149
rect 13181 2964 13211 3164
rect 13432 2970 13462 3194
rect 13976 2968 14006 3192
rect 14079 2968 14109 3168
rect 14180 2989 14210 3189
rect 14281 2947 14311 3147
rect 14371 2947 14401 3147
rect 14468 2947 14498 3147
rect 14585 2947 14615 3147
rect 14686 2947 14716 3147
rect 14778 2947 14808 3147
rect 14879 2947 14909 3147
rect 14969 2947 14999 3147
rect 15088 2947 15118 3147
rect 15255 2962 15285 3162
rect 15506 2968 15536 3192
rect 16038 2964 16068 3188
rect 16141 2964 16171 3164
rect 16242 2985 16272 3185
rect 16343 2943 16373 3143
rect 16433 2943 16463 3143
rect 16530 2943 16560 3143
rect 16647 2943 16677 3143
rect 16748 2943 16778 3143
rect 16840 2943 16870 3143
rect 16941 2943 16971 3143
rect 17031 2943 17061 3143
rect 17150 2943 17180 3143
rect 17317 2958 17347 3158
rect 17568 2964 17598 3188
<< scpmoshvt >>
rect 22664 2883 22694 3083
rect 23249 2881 23279 3081
rect 23333 2881 23363 3081
rect 23865 2869 23895 3069
rect 23949 2869 23979 3069
rect 24033 2869 24063 3069
rect 24117 2869 24147 3069
rect 24713 2855 24743 3055
rect 24797 2855 24827 3055
rect 24881 2855 24911 3055
rect 24965 2855 24995 3055
rect 25049 2855 25079 3055
rect 25133 2855 25163 3055
<< nmoslvt >>
rect 8183 4230 8213 4378
rect 8269 4230 8299 4378
rect 1582 2694 1612 2842
rect 1705 2695 1735 2823
rect 1783 2695 1813 2823
rect 1861 2695 1891 2823
rect 1969 2695 1999 2823
rect 2071 2695 2101 2823
rect 2189 2695 2219 2823
rect 2275 2695 2305 2823
rect 2404 2695 2434 2823
rect 2482 2695 2512 2823
rect 2568 2695 2598 2823
rect 2780 2695 2810 2823
rect 2925 2695 2955 2823
rect 3115 2694 3145 2842
rect 3644 2690 3674 2838
rect 3767 2691 3797 2819
rect 3845 2691 3875 2819
rect 3923 2691 3953 2819
rect 4031 2691 4061 2819
rect 4133 2691 4163 2819
rect 4251 2691 4281 2819
rect 4337 2691 4367 2819
rect 4466 2691 4496 2819
rect 4544 2691 4574 2819
rect 4630 2691 4660 2819
rect 4842 2691 4872 2819
rect 4987 2691 5017 2819
rect 5177 2690 5207 2838
rect 5718 2688 5748 2836
rect 5841 2689 5871 2817
rect 5919 2689 5949 2817
rect 5997 2689 6027 2817
rect 6105 2689 6135 2817
rect 6207 2689 6237 2817
rect 6325 2689 6355 2817
rect 6411 2689 6441 2817
rect 6540 2689 6570 2817
rect 6618 2689 6648 2817
rect 6704 2689 6734 2817
rect 6916 2689 6946 2817
rect 7061 2689 7091 2817
rect 7251 2688 7281 2836
rect 7780 2684 7810 2832
rect 7903 2685 7933 2813
rect 7981 2685 8011 2813
rect 8059 2685 8089 2813
rect 8167 2685 8197 2813
rect 8269 2685 8299 2813
rect 8387 2685 8417 2813
rect 8473 2685 8503 2813
rect 8602 2685 8632 2813
rect 8680 2685 8710 2813
rect 8766 2685 8796 2813
rect 8978 2685 9008 2813
rect 9123 2685 9153 2813
rect 9313 2684 9343 2832
rect 9840 2680 9870 2828
rect 9963 2681 9993 2809
rect 10041 2681 10071 2809
rect 10119 2681 10149 2809
rect 10227 2681 10257 2809
rect 10329 2681 10359 2809
rect 10447 2681 10477 2809
rect 10533 2681 10563 2809
rect 10662 2681 10692 2809
rect 10740 2681 10770 2809
rect 10826 2681 10856 2809
rect 11038 2681 11068 2809
rect 11183 2681 11213 2809
rect 11373 2680 11403 2828
rect 11902 2676 11932 2824
rect 12025 2677 12055 2805
rect 12103 2677 12133 2805
rect 12181 2677 12211 2805
rect 12289 2677 12319 2805
rect 12391 2677 12421 2805
rect 12509 2677 12539 2805
rect 12595 2677 12625 2805
rect 12724 2677 12754 2805
rect 12802 2677 12832 2805
rect 12888 2677 12918 2805
rect 13100 2677 13130 2805
rect 13245 2677 13275 2805
rect 13435 2676 13465 2824
rect 13976 2674 14006 2822
rect 14099 2675 14129 2803
rect 14177 2675 14207 2803
rect 14255 2675 14285 2803
rect 14363 2675 14393 2803
rect 14465 2675 14495 2803
rect 14583 2675 14613 2803
rect 14669 2675 14699 2803
rect 14798 2675 14828 2803
rect 14876 2675 14906 2803
rect 14962 2675 14992 2803
rect 15174 2675 15204 2803
rect 15319 2675 15349 2803
rect 15509 2674 15539 2822
rect 16038 2670 16068 2818
rect 16161 2671 16191 2799
rect 16239 2671 16269 2799
rect 16317 2671 16347 2799
rect 16425 2671 16455 2799
rect 16527 2671 16557 2799
rect 16645 2671 16675 2799
rect 16731 2671 16761 2799
rect 16860 2671 16890 2799
rect 16938 2671 16968 2799
rect 17024 2671 17054 2799
rect 17236 2671 17266 2799
rect 17381 2671 17411 2799
rect 17571 2670 17601 2818
<< ndiff >>
rect 8126 4366 8183 4378
rect 8126 4332 8138 4366
rect 8172 4332 8183 4366
rect 8126 4276 8183 4332
rect 8126 4242 8138 4276
rect 8172 4242 8183 4276
rect 8126 4230 8183 4242
rect 8213 4366 8269 4378
rect 8213 4332 8224 4366
rect 8258 4332 8269 4366
rect 8213 4276 8269 4332
rect 8213 4242 8224 4276
rect 8258 4242 8269 4276
rect 8213 4230 8269 4242
rect 8299 4366 8356 4378
rect 8299 4332 8310 4366
rect 8344 4332 8356 4366
rect 8299 4276 8356 4332
rect 8299 4242 8310 4276
rect 8344 4242 8356 4276
rect 8299 4230 8356 4242
rect 1525 2830 1582 2842
rect 1525 2796 1537 2830
rect 1571 2796 1582 2830
rect 1525 2740 1582 2796
rect 1525 2706 1537 2740
rect 1571 2706 1582 2740
rect 1525 2694 1582 2706
rect 1612 2823 1662 2842
rect 1612 2702 1705 2823
rect 1612 2694 1641 2702
rect 1627 2668 1641 2694
rect 1675 2695 1705 2702
rect 1735 2695 1783 2823
rect 1813 2695 1861 2823
rect 1891 2747 1969 2823
rect 1891 2713 1902 2747
rect 1936 2713 1969 2747
rect 1891 2695 1969 2713
rect 1999 2754 2071 2823
rect 1999 2720 2018 2754
rect 2052 2720 2071 2754
rect 1999 2695 2071 2720
rect 2101 2702 2189 2823
rect 2101 2695 2128 2702
rect 1675 2668 1690 2695
rect 1627 2656 1690 2668
rect 2116 2668 2128 2695
rect 2162 2695 2189 2702
rect 2219 2754 2275 2823
rect 2219 2720 2230 2754
rect 2264 2720 2275 2754
rect 2219 2695 2275 2720
rect 2305 2746 2404 2823
rect 2305 2712 2344 2746
rect 2378 2712 2404 2746
rect 2305 2695 2404 2712
rect 2434 2695 2482 2823
rect 2512 2757 2568 2823
rect 2512 2723 2523 2757
rect 2557 2723 2568 2757
rect 2512 2695 2568 2723
rect 2598 2705 2780 2823
rect 2598 2695 2625 2705
rect 2162 2668 2174 2695
rect 2613 2671 2625 2695
rect 2659 2671 2719 2705
rect 2753 2695 2780 2705
rect 2810 2698 2925 2823
rect 2810 2695 2864 2698
rect 2753 2671 2765 2695
rect 2116 2656 2174 2668
rect 2613 2659 2765 2671
rect 2852 2664 2864 2695
rect 2898 2695 2925 2698
rect 2955 2766 3008 2823
rect 2955 2732 2966 2766
rect 3000 2732 3008 2766
rect 2955 2695 3008 2732
rect 3062 2758 3115 2842
rect 3062 2724 3070 2758
rect 3104 2724 3115 2758
rect 2898 2664 2910 2695
rect 3062 2694 3115 2724
rect 3145 2830 3199 2842
rect 3145 2796 3156 2830
rect 3190 2796 3199 2830
rect 3145 2740 3199 2796
rect 3145 2706 3156 2740
rect 3190 2706 3199 2740
rect 3145 2694 3199 2706
rect 3587 2826 3644 2838
rect 3587 2792 3599 2826
rect 3633 2792 3644 2826
rect 3587 2736 3644 2792
rect 3587 2702 3599 2736
rect 3633 2702 3644 2736
rect 3587 2690 3644 2702
rect 3674 2819 3724 2838
rect 3674 2698 3767 2819
rect 3674 2690 3703 2698
rect 3689 2664 3703 2690
rect 3737 2691 3767 2698
rect 3797 2691 3845 2819
rect 3875 2691 3923 2819
rect 3953 2743 4031 2819
rect 3953 2709 3964 2743
rect 3998 2709 4031 2743
rect 3953 2691 4031 2709
rect 4061 2750 4133 2819
rect 4061 2716 4080 2750
rect 4114 2716 4133 2750
rect 4061 2691 4133 2716
rect 4163 2698 4251 2819
rect 4163 2691 4190 2698
rect 3737 2664 3752 2691
rect 2852 2656 2910 2664
rect 3689 2652 3752 2664
rect 4178 2664 4190 2691
rect 4224 2691 4251 2698
rect 4281 2750 4337 2819
rect 4281 2716 4292 2750
rect 4326 2716 4337 2750
rect 4281 2691 4337 2716
rect 4367 2742 4466 2819
rect 4367 2708 4406 2742
rect 4440 2708 4466 2742
rect 4367 2691 4466 2708
rect 4496 2691 4544 2819
rect 4574 2753 4630 2819
rect 4574 2719 4585 2753
rect 4619 2719 4630 2753
rect 4574 2691 4630 2719
rect 4660 2701 4842 2819
rect 4660 2691 4687 2701
rect 4224 2664 4236 2691
rect 4675 2667 4687 2691
rect 4721 2667 4781 2701
rect 4815 2691 4842 2701
rect 4872 2694 4987 2819
rect 4872 2691 4926 2694
rect 4815 2667 4827 2691
rect 4178 2652 4236 2664
rect 4675 2655 4827 2667
rect 4914 2660 4926 2691
rect 4960 2691 4987 2694
rect 5017 2762 5070 2819
rect 5017 2728 5028 2762
rect 5062 2728 5070 2762
rect 5017 2691 5070 2728
rect 5124 2754 5177 2838
rect 5124 2720 5132 2754
rect 5166 2720 5177 2754
rect 4960 2660 4972 2691
rect 5124 2690 5177 2720
rect 5207 2826 5261 2838
rect 5207 2792 5218 2826
rect 5252 2792 5261 2826
rect 5207 2736 5261 2792
rect 5207 2702 5218 2736
rect 5252 2702 5261 2736
rect 5207 2690 5261 2702
rect 5661 2824 5718 2836
rect 5661 2790 5673 2824
rect 5707 2790 5718 2824
rect 5661 2734 5718 2790
rect 5661 2700 5673 2734
rect 5707 2700 5718 2734
rect 5661 2688 5718 2700
rect 5748 2817 5798 2836
rect 5748 2696 5841 2817
rect 5748 2688 5777 2696
rect 5763 2662 5777 2688
rect 5811 2689 5841 2696
rect 5871 2689 5919 2817
rect 5949 2689 5997 2817
rect 6027 2741 6105 2817
rect 6027 2707 6038 2741
rect 6072 2707 6105 2741
rect 6027 2689 6105 2707
rect 6135 2748 6207 2817
rect 6135 2714 6154 2748
rect 6188 2714 6207 2748
rect 6135 2689 6207 2714
rect 6237 2696 6325 2817
rect 6237 2689 6264 2696
rect 5811 2662 5826 2689
rect 4914 2652 4972 2660
rect 5763 2650 5826 2662
rect 6252 2662 6264 2689
rect 6298 2689 6325 2696
rect 6355 2748 6411 2817
rect 6355 2714 6366 2748
rect 6400 2714 6411 2748
rect 6355 2689 6411 2714
rect 6441 2740 6540 2817
rect 6441 2706 6480 2740
rect 6514 2706 6540 2740
rect 6441 2689 6540 2706
rect 6570 2689 6618 2817
rect 6648 2751 6704 2817
rect 6648 2717 6659 2751
rect 6693 2717 6704 2751
rect 6648 2689 6704 2717
rect 6734 2699 6916 2817
rect 6734 2689 6761 2699
rect 6298 2662 6310 2689
rect 6749 2665 6761 2689
rect 6795 2665 6855 2699
rect 6889 2689 6916 2699
rect 6946 2692 7061 2817
rect 6946 2689 7000 2692
rect 6889 2665 6901 2689
rect 6252 2650 6310 2662
rect 6749 2653 6901 2665
rect 6988 2658 7000 2689
rect 7034 2689 7061 2692
rect 7091 2760 7144 2817
rect 7091 2726 7102 2760
rect 7136 2726 7144 2760
rect 7091 2689 7144 2726
rect 7198 2752 7251 2836
rect 7198 2718 7206 2752
rect 7240 2718 7251 2752
rect 7034 2658 7046 2689
rect 7198 2688 7251 2718
rect 7281 2824 7335 2836
rect 7281 2790 7292 2824
rect 7326 2790 7335 2824
rect 7281 2734 7335 2790
rect 7281 2700 7292 2734
rect 7326 2700 7335 2734
rect 7281 2688 7335 2700
rect 7723 2820 7780 2832
rect 7723 2786 7735 2820
rect 7769 2786 7780 2820
rect 7723 2730 7780 2786
rect 7723 2696 7735 2730
rect 7769 2696 7780 2730
rect 7723 2684 7780 2696
rect 7810 2813 7860 2832
rect 7810 2692 7903 2813
rect 7810 2684 7839 2692
rect 7825 2658 7839 2684
rect 7873 2685 7903 2692
rect 7933 2685 7981 2813
rect 8011 2685 8059 2813
rect 8089 2737 8167 2813
rect 8089 2703 8100 2737
rect 8134 2703 8167 2737
rect 8089 2685 8167 2703
rect 8197 2744 8269 2813
rect 8197 2710 8216 2744
rect 8250 2710 8269 2744
rect 8197 2685 8269 2710
rect 8299 2692 8387 2813
rect 8299 2685 8326 2692
rect 7873 2658 7888 2685
rect 6988 2650 7046 2658
rect 7825 2646 7888 2658
rect 8314 2658 8326 2685
rect 8360 2685 8387 2692
rect 8417 2744 8473 2813
rect 8417 2710 8428 2744
rect 8462 2710 8473 2744
rect 8417 2685 8473 2710
rect 8503 2736 8602 2813
rect 8503 2702 8542 2736
rect 8576 2702 8602 2736
rect 8503 2685 8602 2702
rect 8632 2685 8680 2813
rect 8710 2747 8766 2813
rect 8710 2713 8721 2747
rect 8755 2713 8766 2747
rect 8710 2685 8766 2713
rect 8796 2695 8978 2813
rect 8796 2685 8823 2695
rect 8360 2658 8372 2685
rect 8811 2661 8823 2685
rect 8857 2661 8917 2695
rect 8951 2685 8978 2695
rect 9008 2688 9123 2813
rect 9008 2685 9062 2688
rect 8951 2661 8963 2685
rect 8314 2646 8372 2658
rect 8811 2649 8963 2661
rect 9050 2654 9062 2685
rect 9096 2685 9123 2688
rect 9153 2756 9206 2813
rect 9153 2722 9164 2756
rect 9198 2722 9206 2756
rect 9153 2685 9206 2722
rect 9260 2748 9313 2832
rect 9260 2714 9268 2748
rect 9302 2714 9313 2748
rect 9096 2654 9108 2685
rect 9260 2684 9313 2714
rect 9343 2820 9397 2832
rect 9343 2786 9354 2820
rect 9388 2786 9397 2820
rect 9343 2730 9397 2786
rect 9343 2696 9354 2730
rect 9388 2696 9397 2730
rect 9343 2684 9397 2696
rect 9783 2816 9840 2828
rect 9783 2782 9795 2816
rect 9829 2782 9840 2816
rect 9783 2726 9840 2782
rect 9783 2692 9795 2726
rect 9829 2692 9840 2726
rect 9783 2680 9840 2692
rect 9870 2809 9920 2828
rect 9870 2688 9963 2809
rect 9870 2680 9899 2688
rect 9885 2654 9899 2680
rect 9933 2681 9963 2688
rect 9993 2681 10041 2809
rect 10071 2681 10119 2809
rect 10149 2733 10227 2809
rect 10149 2699 10160 2733
rect 10194 2699 10227 2733
rect 10149 2681 10227 2699
rect 10257 2740 10329 2809
rect 10257 2706 10276 2740
rect 10310 2706 10329 2740
rect 10257 2681 10329 2706
rect 10359 2688 10447 2809
rect 10359 2681 10386 2688
rect 9933 2654 9948 2681
rect 9050 2646 9108 2654
rect 9885 2642 9948 2654
rect 10374 2654 10386 2681
rect 10420 2681 10447 2688
rect 10477 2740 10533 2809
rect 10477 2706 10488 2740
rect 10522 2706 10533 2740
rect 10477 2681 10533 2706
rect 10563 2732 10662 2809
rect 10563 2698 10602 2732
rect 10636 2698 10662 2732
rect 10563 2681 10662 2698
rect 10692 2681 10740 2809
rect 10770 2743 10826 2809
rect 10770 2709 10781 2743
rect 10815 2709 10826 2743
rect 10770 2681 10826 2709
rect 10856 2691 11038 2809
rect 10856 2681 10883 2691
rect 10420 2654 10432 2681
rect 10871 2657 10883 2681
rect 10917 2657 10977 2691
rect 11011 2681 11038 2691
rect 11068 2684 11183 2809
rect 11068 2681 11122 2684
rect 11011 2657 11023 2681
rect 10374 2642 10432 2654
rect 10871 2645 11023 2657
rect 11110 2650 11122 2681
rect 11156 2681 11183 2684
rect 11213 2752 11266 2809
rect 11213 2718 11224 2752
rect 11258 2718 11266 2752
rect 11213 2681 11266 2718
rect 11320 2744 11373 2828
rect 11320 2710 11328 2744
rect 11362 2710 11373 2744
rect 11156 2650 11168 2681
rect 11320 2680 11373 2710
rect 11403 2816 11457 2828
rect 11403 2782 11414 2816
rect 11448 2782 11457 2816
rect 11403 2726 11457 2782
rect 11403 2692 11414 2726
rect 11448 2692 11457 2726
rect 11403 2680 11457 2692
rect 11845 2812 11902 2824
rect 11845 2778 11857 2812
rect 11891 2778 11902 2812
rect 11845 2722 11902 2778
rect 11845 2688 11857 2722
rect 11891 2688 11902 2722
rect 11845 2676 11902 2688
rect 11932 2805 11982 2824
rect 11932 2684 12025 2805
rect 11932 2676 11961 2684
rect 11947 2650 11961 2676
rect 11995 2677 12025 2684
rect 12055 2677 12103 2805
rect 12133 2677 12181 2805
rect 12211 2729 12289 2805
rect 12211 2695 12222 2729
rect 12256 2695 12289 2729
rect 12211 2677 12289 2695
rect 12319 2736 12391 2805
rect 12319 2702 12338 2736
rect 12372 2702 12391 2736
rect 12319 2677 12391 2702
rect 12421 2684 12509 2805
rect 12421 2677 12448 2684
rect 11995 2650 12010 2677
rect 11110 2642 11168 2650
rect 11947 2638 12010 2650
rect 12436 2650 12448 2677
rect 12482 2677 12509 2684
rect 12539 2736 12595 2805
rect 12539 2702 12550 2736
rect 12584 2702 12595 2736
rect 12539 2677 12595 2702
rect 12625 2728 12724 2805
rect 12625 2694 12664 2728
rect 12698 2694 12724 2728
rect 12625 2677 12724 2694
rect 12754 2677 12802 2805
rect 12832 2739 12888 2805
rect 12832 2705 12843 2739
rect 12877 2705 12888 2739
rect 12832 2677 12888 2705
rect 12918 2687 13100 2805
rect 12918 2677 12945 2687
rect 12482 2650 12494 2677
rect 12933 2653 12945 2677
rect 12979 2653 13039 2687
rect 13073 2677 13100 2687
rect 13130 2680 13245 2805
rect 13130 2677 13184 2680
rect 13073 2653 13085 2677
rect 12436 2638 12494 2650
rect 12933 2641 13085 2653
rect 13172 2646 13184 2677
rect 13218 2677 13245 2680
rect 13275 2748 13328 2805
rect 13275 2714 13286 2748
rect 13320 2714 13328 2748
rect 13275 2677 13328 2714
rect 13382 2740 13435 2824
rect 13382 2706 13390 2740
rect 13424 2706 13435 2740
rect 13218 2646 13230 2677
rect 13382 2676 13435 2706
rect 13465 2812 13519 2824
rect 13465 2778 13476 2812
rect 13510 2778 13519 2812
rect 13465 2722 13519 2778
rect 13465 2688 13476 2722
rect 13510 2688 13519 2722
rect 13465 2676 13519 2688
rect 13919 2810 13976 2822
rect 13919 2776 13931 2810
rect 13965 2776 13976 2810
rect 13919 2720 13976 2776
rect 13919 2686 13931 2720
rect 13965 2686 13976 2720
rect 13919 2674 13976 2686
rect 14006 2803 14056 2822
rect 14006 2682 14099 2803
rect 14006 2674 14035 2682
rect 14021 2648 14035 2674
rect 14069 2675 14099 2682
rect 14129 2675 14177 2803
rect 14207 2675 14255 2803
rect 14285 2727 14363 2803
rect 14285 2693 14296 2727
rect 14330 2693 14363 2727
rect 14285 2675 14363 2693
rect 14393 2734 14465 2803
rect 14393 2700 14412 2734
rect 14446 2700 14465 2734
rect 14393 2675 14465 2700
rect 14495 2682 14583 2803
rect 14495 2675 14522 2682
rect 14069 2648 14084 2675
rect 13172 2638 13230 2646
rect 14021 2636 14084 2648
rect 14510 2648 14522 2675
rect 14556 2675 14583 2682
rect 14613 2734 14669 2803
rect 14613 2700 14624 2734
rect 14658 2700 14669 2734
rect 14613 2675 14669 2700
rect 14699 2726 14798 2803
rect 14699 2692 14738 2726
rect 14772 2692 14798 2726
rect 14699 2675 14798 2692
rect 14828 2675 14876 2803
rect 14906 2737 14962 2803
rect 14906 2703 14917 2737
rect 14951 2703 14962 2737
rect 14906 2675 14962 2703
rect 14992 2685 15174 2803
rect 14992 2675 15019 2685
rect 14556 2648 14568 2675
rect 15007 2651 15019 2675
rect 15053 2651 15113 2685
rect 15147 2675 15174 2685
rect 15204 2678 15319 2803
rect 15204 2675 15258 2678
rect 15147 2651 15159 2675
rect 14510 2636 14568 2648
rect 15007 2639 15159 2651
rect 15246 2644 15258 2675
rect 15292 2675 15319 2678
rect 15349 2746 15402 2803
rect 15349 2712 15360 2746
rect 15394 2712 15402 2746
rect 15349 2675 15402 2712
rect 15456 2738 15509 2822
rect 15456 2704 15464 2738
rect 15498 2704 15509 2738
rect 15292 2644 15304 2675
rect 15456 2674 15509 2704
rect 15539 2810 15593 2822
rect 15539 2776 15550 2810
rect 15584 2776 15593 2810
rect 15539 2720 15593 2776
rect 15539 2686 15550 2720
rect 15584 2686 15593 2720
rect 15539 2674 15593 2686
rect 15981 2806 16038 2818
rect 15981 2772 15993 2806
rect 16027 2772 16038 2806
rect 15981 2716 16038 2772
rect 15981 2682 15993 2716
rect 16027 2682 16038 2716
rect 15981 2670 16038 2682
rect 16068 2799 16118 2818
rect 16068 2678 16161 2799
rect 16068 2670 16097 2678
rect 16083 2644 16097 2670
rect 16131 2671 16161 2678
rect 16191 2671 16239 2799
rect 16269 2671 16317 2799
rect 16347 2723 16425 2799
rect 16347 2689 16358 2723
rect 16392 2689 16425 2723
rect 16347 2671 16425 2689
rect 16455 2730 16527 2799
rect 16455 2696 16474 2730
rect 16508 2696 16527 2730
rect 16455 2671 16527 2696
rect 16557 2678 16645 2799
rect 16557 2671 16584 2678
rect 16131 2644 16146 2671
rect 15246 2636 15304 2644
rect 16083 2632 16146 2644
rect 16572 2644 16584 2671
rect 16618 2671 16645 2678
rect 16675 2730 16731 2799
rect 16675 2696 16686 2730
rect 16720 2696 16731 2730
rect 16675 2671 16731 2696
rect 16761 2722 16860 2799
rect 16761 2688 16800 2722
rect 16834 2688 16860 2722
rect 16761 2671 16860 2688
rect 16890 2671 16938 2799
rect 16968 2733 17024 2799
rect 16968 2699 16979 2733
rect 17013 2699 17024 2733
rect 16968 2671 17024 2699
rect 17054 2681 17236 2799
rect 17054 2671 17081 2681
rect 16618 2644 16630 2671
rect 17069 2647 17081 2671
rect 17115 2647 17175 2681
rect 17209 2671 17236 2681
rect 17266 2674 17381 2799
rect 17266 2671 17320 2674
rect 17209 2647 17221 2671
rect 16572 2632 16630 2644
rect 17069 2635 17221 2647
rect 17308 2640 17320 2671
rect 17354 2671 17381 2674
rect 17411 2742 17464 2799
rect 17411 2708 17422 2742
rect 17456 2708 17464 2742
rect 17411 2671 17464 2708
rect 17518 2734 17571 2818
rect 17518 2700 17526 2734
rect 17560 2700 17571 2734
rect 17354 2640 17366 2671
rect 17518 2670 17571 2700
rect 17601 2806 17655 2818
rect 17601 2772 17612 2806
rect 17646 2772 17655 2806
rect 17601 2716 17655 2772
rect 17601 2682 17612 2716
rect 17646 2682 17655 2716
rect 17601 2670 17655 2682
rect 22612 2751 22664 2763
rect 22612 2717 22620 2751
rect 22654 2717 22664 2751
rect 22612 2683 22664 2717
rect 22612 2649 22620 2683
rect 22654 2649 22664 2683
rect 17308 2632 17366 2640
rect 22612 2633 22664 2649
rect 22694 2751 22746 2763
rect 22694 2717 22704 2751
rect 22738 2717 22746 2751
rect 22694 2683 22746 2717
rect 22694 2649 22704 2683
rect 22738 2649 22746 2683
rect 22694 2633 22746 2649
rect 23197 2749 23249 2761
rect 23197 2715 23205 2749
rect 23239 2715 23249 2749
rect 23197 2677 23249 2715
rect 23197 2643 23205 2677
rect 23239 2643 23249 2677
rect 23197 2631 23249 2643
rect 23279 2749 23333 2761
rect 23279 2715 23289 2749
rect 23323 2715 23333 2749
rect 23279 2677 23333 2715
rect 23279 2643 23289 2677
rect 23323 2643 23333 2677
rect 23279 2631 23333 2643
rect 23363 2749 23415 2761
rect 23363 2715 23373 2749
rect 23407 2715 23415 2749
rect 23363 2677 23415 2715
rect 23363 2643 23373 2677
rect 23407 2643 23415 2677
rect 23363 2631 23415 2643
rect 23813 2665 23865 2749
rect 23813 2631 23821 2665
rect 23855 2631 23865 2665
rect 23813 2619 23865 2631
rect 23895 2673 23949 2749
rect 23895 2639 23905 2673
rect 23939 2639 23949 2673
rect 23895 2619 23949 2639
rect 23979 2665 24033 2749
rect 23979 2631 23989 2665
rect 24023 2631 24033 2665
rect 23979 2619 24033 2631
rect 24063 2673 24117 2749
rect 24063 2639 24073 2673
rect 24107 2639 24117 2673
rect 24063 2619 24117 2639
rect 24147 2666 24199 2749
rect 24147 2632 24157 2666
rect 24191 2632 24199 2666
rect 24147 2619 24199 2632
rect 24637 2651 24713 2735
rect 24637 2617 24645 2651
rect 24679 2617 24713 2651
rect 24637 2605 24713 2617
rect 24743 2659 24797 2735
rect 24743 2625 24753 2659
rect 24787 2625 24797 2659
rect 24743 2605 24797 2625
rect 24827 2651 24881 2735
rect 24827 2617 24837 2651
rect 24871 2617 24881 2651
rect 24827 2605 24881 2617
rect 24911 2659 24965 2735
rect 24911 2625 24921 2659
rect 24955 2625 24965 2659
rect 24911 2605 24965 2625
rect 24995 2651 25049 2735
rect 24995 2617 25005 2651
rect 25039 2617 25049 2651
rect 24995 2605 25049 2617
rect 25079 2659 25133 2735
rect 25079 2625 25089 2659
rect 25123 2625 25133 2659
rect 25079 2605 25133 2625
rect 25163 2652 25217 2735
rect 25163 2618 25173 2652
rect 25207 2618 25217 2652
rect 25163 2605 25217 2618
<< pdiff >>
rect 8125 4072 8182 4084
rect 8125 4038 8135 4072
rect 8169 4038 8182 4072
rect 8125 3989 8182 4038
rect 8125 3955 8135 3989
rect 8169 3955 8182 3989
rect 8125 3906 8182 3955
rect 8125 3872 8135 3906
rect 8169 3872 8182 3906
rect 8125 3860 8182 3872
rect 8212 4072 8272 4084
rect 8212 4038 8225 4072
rect 8259 4038 8272 4072
rect 8212 3989 8272 4038
rect 8212 3955 8225 3989
rect 8259 3955 8272 3989
rect 8212 3906 8272 3955
rect 8212 3872 8225 3906
rect 8259 3872 8272 3906
rect 8212 3860 8272 3872
rect 8302 4046 8359 4084
rect 8302 4012 8315 4046
rect 8349 4012 8359 4046
rect 8302 3976 8359 4012
rect 8302 3942 8315 3976
rect 8349 3942 8359 3976
rect 8302 3906 8359 3942
rect 8302 3872 8315 3906
rect 8349 3872 8359 3906
rect 8302 3860 8359 3872
rect 1525 3200 1582 3212
rect 1525 3166 1535 3200
rect 1569 3166 1582 3200
rect 1525 3117 1582 3166
rect 1525 3083 1535 3117
rect 1569 3083 1582 3117
rect 1525 3034 1582 3083
rect 1525 3000 1535 3034
rect 1569 3000 1582 3034
rect 1525 2988 1582 3000
rect 1612 3200 1667 3212
rect 1612 3166 1625 3200
rect 1659 3188 1667 3200
rect 1733 3188 1786 3209
rect 1659 3166 1685 3188
rect 1612 3132 1685 3166
rect 1612 3098 1625 3132
rect 1659 3098 1685 3132
rect 1612 3064 1685 3098
rect 1612 3030 1625 3064
rect 1659 3030 1685 3064
rect 1612 2988 1685 3030
rect 1715 3009 1786 3188
rect 1816 3167 1869 3209
rect 2122 3196 2173 3208
rect 2122 3167 2130 3196
rect 1816 3009 1887 3167
rect 1715 2988 1768 3009
rect 1834 2967 1887 3009
rect 1917 3155 1977 3167
rect 1917 3121 1930 3155
rect 1964 3121 1977 3155
rect 1917 3087 1977 3121
rect 1917 3053 1930 3087
rect 1964 3053 1977 3087
rect 1917 3019 1977 3053
rect 1917 2985 1930 3019
rect 1964 2985 1977 3019
rect 1917 2967 1977 2985
rect 2007 3155 2074 3167
rect 2007 3121 2020 3155
rect 2054 3121 2074 3155
rect 2007 3063 2074 3121
rect 2007 3029 2020 3063
rect 2054 3029 2074 3063
rect 2007 2967 2074 3029
rect 2104 3162 2130 3167
rect 2164 3167 2173 3196
rect 3053 3200 3112 3212
rect 2742 3167 2861 3182
rect 2164 3162 2191 3167
rect 2104 2967 2191 3162
rect 2221 3128 2292 3167
rect 2221 3094 2234 3128
rect 2268 3094 2292 3128
rect 2221 2967 2292 3094
rect 2322 3131 2384 3167
rect 2322 3097 2335 3131
rect 2369 3097 2384 3131
rect 2322 2967 2384 3097
rect 2414 2967 2485 3167
rect 2515 3155 2575 3167
rect 2515 3121 2528 3155
rect 2562 3121 2575 3155
rect 2515 3044 2575 3121
rect 2515 3010 2528 3044
rect 2562 3010 2575 3044
rect 2515 2967 2575 3010
rect 2605 3155 2694 3167
rect 2605 3121 2647 3155
rect 2681 3121 2694 3155
rect 2605 3071 2694 3121
rect 2605 3037 2647 3071
rect 2681 3037 2694 3071
rect 2605 2967 2694 3037
rect 2724 3157 2861 3167
rect 2724 3123 2738 3157
rect 2772 3123 2813 3157
rect 2847 3123 2861 3157
rect 2724 2982 2861 3123
rect 2891 3170 2958 3182
rect 2891 3136 2912 3170
rect 2946 3136 2958 3170
rect 2891 3060 2958 3136
rect 2891 3026 2912 3060
rect 2946 3026 2958 3060
rect 2891 2982 2958 3026
rect 3053 3166 3065 3200
rect 3099 3166 3112 3200
rect 3053 3117 3112 3166
rect 3053 3083 3065 3117
rect 3099 3083 3112 3117
rect 3053 3034 3112 3083
rect 3053 3000 3065 3034
rect 3099 3000 3112 3034
rect 3053 2988 3112 3000
rect 3142 3200 3199 3212
rect 3142 3166 3155 3200
rect 3189 3166 3199 3200
rect 3142 3117 3199 3166
rect 3142 3083 3155 3117
rect 3189 3083 3199 3117
rect 3142 3034 3199 3083
rect 3142 3000 3155 3034
rect 3189 3000 3199 3034
rect 3142 2988 3199 3000
rect 3587 3196 3644 3208
rect 3587 3162 3597 3196
rect 3631 3162 3644 3196
rect 3587 3113 3644 3162
rect 3587 3079 3597 3113
rect 3631 3079 3644 3113
rect 3587 3030 3644 3079
rect 3587 2996 3597 3030
rect 3631 2996 3644 3030
rect 2724 2967 2777 2982
rect 3587 2984 3644 2996
rect 3674 3196 3729 3208
rect 3674 3162 3687 3196
rect 3721 3184 3729 3196
rect 3795 3184 3848 3205
rect 3721 3162 3747 3184
rect 3674 3128 3747 3162
rect 3674 3094 3687 3128
rect 3721 3094 3747 3128
rect 3674 3060 3747 3094
rect 3674 3026 3687 3060
rect 3721 3026 3747 3060
rect 3674 2984 3747 3026
rect 3777 3005 3848 3184
rect 3878 3163 3931 3205
rect 4184 3192 4235 3204
rect 4184 3163 4192 3192
rect 3878 3005 3949 3163
rect 3777 2984 3830 3005
rect 3896 2963 3949 3005
rect 3979 3151 4039 3163
rect 3979 3117 3992 3151
rect 4026 3117 4039 3151
rect 3979 3083 4039 3117
rect 3979 3049 3992 3083
rect 4026 3049 4039 3083
rect 3979 3015 4039 3049
rect 3979 2981 3992 3015
rect 4026 2981 4039 3015
rect 3979 2963 4039 2981
rect 4069 3151 4136 3163
rect 4069 3117 4082 3151
rect 4116 3117 4136 3151
rect 4069 3059 4136 3117
rect 4069 3025 4082 3059
rect 4116 3025 4136 3059
rect 4069 2963 4136 3025
rect 4166 3158 4192 3163
rect 4226 3163 4235 3192
rect 5115 3196 5174 3208
rect 4804 3163 4923 3178
rect 4226 3158 4253 3163
rect 4166 2963 4253 3158
rect 4283 3124 4354 3163
rect 4283 3090 4296 3124
rect 4330 3090 4354 3124
rect 4283 2963 4354 3090
rect 4384 3127 4446 3163
rect 4384 3093 4397 3127
rect 4431 3093 4446 3127
rect 4384 2963 4446 3093
rect 4476 2963 4547 3163
rect 4577 3151 4637 3163
rect 4577 3117 4590 3151
rect 4624 3117 4637 3151
rect 4577 3040 4637 3117
rect 4577 3006 4590 3040
rect 4624 3006 4637 3040
rect 4577 2963 4637 3006
rect 4667 3151 4756 3163
rect 4667 3117 4709 3151
rect 4743 3117 4756 3151
rect 4667 3067 4756 3117
rect 4667 3033 4709 3067
rect 4743 3033 4756 3067
rect 4667 2963 4756 3033
rect 4786 3153 4923 3163
rect 4786 3119 4800 3153
rect 4834 3119 4875 3153
rect 4909 3119 4923 3153
rect 4786 2978 4923 3119
rect 4953 3166 5020 3178
rect 4953 3132 4974 3166
rect 5008 3132 5020 3166
rect 4953 3056 5020 3132
rect 4953 3022 4974 3056
rect 5008 3022 5020 3056
rect 4953 2978 5020 3022
rect 5115 3162 5127 3196
rect 5161 3162 5174 3196
rect 5115 3113 5174 3162
rect 5115 3079 5127 3113
rect 5161 3079 5174 3113
rect 5115 3030 5174 3079
rect 5115 2996 5127 3030
rect 5161 2996 5174 3030
rect 5115 2984 5174 2996
rect 5204 3196 5261 3208
rect 5204 3162 5217 3196
rect 5251 3162 5261 3196
rect 5204 3113 5261 3162
rect 5204 3079 5217 3113
rect 5251 3079 5261 3113
rect 5204 3030 5261 3079
rect 5204 2996 5217 3030
rect 5251 2996 5261 3030
rect 5204 2984 5261 2996
rect 5661 3194 5718 3206
rect 5661 3160 5671 3194
rect 5705 3160 5718 3194
rect 5661 3111 5718 3160
rect 5661 3077 5671 3111
rect 5705 3077 5718 3111
rect 5661 3028 5718 3077
rect 5661 2994 5671 3028
rect 5705 2994 5718 3028
rect 4786 2963 4839 2978
rect 5661 2982 5718 2994
rect 5748 3194 5803 3206
rect 5748 3160 5761 3194
rect 5795 3182 5803 3194
rect 5869 3182 5922 3203
rect 5795 3160 5821 3182
rect 5748 3126 5821 3160
rect 5748 3092 5761 3126
rect 5795 3092 5821 3126
rect 5748 3058 5821 3092
rect 5748 3024 5761 3058
rect 5795 3024 5821 3058
rect 5748 2982 5821 3024
rect 5851 3003 5922 3182
rect 5952 3161 6005 3203
rect 6258 3190 6309 3202
rect 6258 3161 6266 3190
rect 5952 3003 6023 3161
rect 5851 2982 5904 3003
rect 5970 2961 6023 3003
rect 6053 3149 6113 3161
rect 6053 3115 6066 3149
rect 6100 3115 6113 3149
rect 6053 3081 6113 3115
rect 6053 3047 6066 3081
rect 6100 3047 6113 3081
rect 6053 3013 6113 3047
rect 6053 2979 6066 3013
rect 6100 2979 6113 3013
rect 6053 2961 6113 2979
rect 6143 3149 6210 3161
rect 6143 3115 6156 3149
rect 6190 3115 6210 3149
rect 6143 3057 6210 3115
rect 6143 3023 6156 3057
rect 6190 3023 6210 3057
rect 6143 2961 6210 3023
rect 6240 3156 6266 3161
rect 6300 3161 6309 3190
rect 7189 3194 7248 3206
rect 6878 3161 6997 3176
rect 6300 3156 6327 3161
rect 6240 2961 6327 3156
rect 6357 3122 6428 3161
rect 6357 3088 6370 3122
rect 6404 3088 6428 3122
rect 6357 2961 6428 3088
rect 6458 3125 6520 3161
rect 6458 3091 6471 3125
rect 6505 3091 6520 3125
rect 6458 2961 6520 3091
rect 6550 2961 6621 3161
rect 6651 3149 6711 3161
rect 6651 3115 6664 3149
rect 6698 3115 6711 3149
rect 6651 3038 6711 3115
rect 6651 3004 6664 3038
rect 6698 3004 6711 3038
rect 6651 2961 6711 3004
rect 6741 3149 6830 3161
rect 6741 3115 6783 3149
rect 6817 3115 6830 3149
rect 6741 3065 6830 3115
rect 6741 3031 6783 3065
rect 6817 3031 6830 3065
rect 6741 2961 6830 3031
rect 6860 3151 6997 3161
rect 6860 3117 6874 3151
rect 6908 3117 6949 3151
rect 6983 3117 6997 3151
rect 6860 2976 6997 3117
rect 7027 3164 7094 3176
rect 7027 3130 7048 3164
rect 7082 3130 7094 3164
rect 7027 3054 7094 3130
rect 7027 3020 7048 3054
rect 7082 3020 7094 3054
rect 7027 2976 7094 3020
rect 7189 3160 7201 3194
rect 7235 3160 7248 3194
rect 7189 3111 7248 3160
rect 7189 3077 7201 3111
rect 7235 3077 7248 3111
rect 7189 3028 7248 3077
rect 7189 2994 7201 3028
rect 7235 2994 7248 3028
rect 7189 2982 7248 2994
rect 7278 3194 7335 3206
rect 7278 3160 7291 3194
rect 7325 3160 7335 3194
rect 7278 3111 7335 3160
rect 7278 3077 7291 3111
rect 7325 3077 7335 3111
rect 7278 3028 7335 3077
rect 7278 2994 7291 3028
rect 7325 2994 7335 3028
rect 7278 2982 7335 2994
rect 7723 3190 7780 3202
rect 7723 3156 7733 3190
rect 7767 3156 7780 3190
rect 7723 3107 7780 3156
rect 7723 3073 7733 3107
rect 7767 3073 7780 3107
rect 7723 3024 7780 3073
rect 7723 2990 7733 3024
rect 7767 2990 7780 3024
rect 6860 2961 6913 2976
rect 7723 2978 7780 2990
rect 7810 3190 7865 3202
rect 7810 3156 7823 3190
rect 7857 3178 7865 3190
rect 7931 3178 7984 3199
rect 7857 3156 7883 3178
rect 7810 3122 7883 3156
rect 7810 3088 7823 3122
rect 7857 3088 7883 3122
rect 7810 3054 7883 3088
rect 7810 3020 7823 3054
rect 7857 3020 7883 3054
rect 7810 2978 7883 3020
rect 7913 2999 7984 3178
rect 8014 3157 8067 3199
rect 8320 3186 8371 3198
rect 8320 3157 8328 3186
rect 8014 2999 8085 3157
rect 7913 2978 7966 2999
rect 8032 2957 8085 2999
rect 8115 3145 8175 3157
rect 8115 3111 8128 3145
rect 8162 3111 8175 3145
rect 8115 3077 8175 3111
rect 8115 3043 8128 3077
rect 8162 3043 8175 3077
rect 8115 3009 8175 3043
rect 8115 2975 8128 3009
rect 8162 2975 8175 3009
rect 8115 2957 8175 2975
rect 8205 3145 8272 3157
rect 8205 3111 8218 3145
rect 8252 3111 8272 3145
rect 8205 3053 8272 3111
rect 8205 3019 8218 3053
rect 8252 3019 8272 3053
rect 8205 2957 8272 3019
rect 8302 3152 8328 3157
rect 8362 3157 8371 3186
rect 9251 3190 9310 3202
rect 8940 3157 9059 3172
rect 8362 3152 8389 3157
rect 8302 2957 8389 3152
rect 8419 3118 8490 3157
rect 8419 3084 8432 3118
rect 8466 3084 8490 3118
rect 8419 2957 8490 3084
rect 8520 3121 8582 3157
rect 8520 3087 8533 3121
rect 8567 3087 8582 3121
rect 8520 2957 8582 3087
rect 8612 2957 8683 3157
rect 8713 3145 8773 3157
rect 8713 3111 8726 3145
rect 8760 3111 8773 3145
rect 8713 3034 8773 3111
rect 8713 3000 8726 3034
rect 8760 3000 8773 3034
rect 8713 2957 8773 3000
rect 8803 3145 8892 3157
rect 8803 3111 8845 3145
rect 8879 3111 8892 3145
rect 8803 3061 8892 3111
rect 8803 3027 8845 3061
rect 8879 3027 8892 3061
rect 8803 2957 8892 3027
rect 8922 3147 9059 3157
rect 8922 3113 8936 3147
rect 8970 3113 9011 3147
rect 9045 3113 9059 3147
rect 8922 2972 9059 3113
rect 9089 3160 9156 3172
rect 9089 3126 9110 3160
rect 9144 3126 9156 3160
rect 9089 3050 9156 3126
rect 9089 3016 9110 3050
rect 9144 3016 9156 3050
rect 9089 2972 9156 3016
rect 9251 3156 9263 3190
rect 9297 3156 9310 3190
rect 9251 3107 9310 3156
rect 9251 3073 9263 3107
rect 9297 3073 9310 3107
rect 9251 3024 9310 3073
rect 9251 2990 9263 3024
rect 9297 2990 9310 3024
rect 9251 2978 9310 2990
rect 9340 3190 9397 3202
rect 9340 3156 9353 3190
rect 9387 3156 9397 3190
rect 9340 3107 9397 3156
rect 9340 3073 9353 3107
rect 9387 3073 9397 3107
rect 9340 3024 9397 3073
rect 9340 2990 9353 3024
rect 9387 2990 9397 3024
rect 9340 2978 9397 2990
rect 9783 3186 9840 3198
rect 9783 3152 9793 3186
rect 9827 3152 9840 3186
rect 9783 3103 9840 3152
rect 9783 3069 9793 3103
rect 9827 3069 9840 3103
rect 9783 3020 9840 3069
rect 9783 2986 9793 3020
rect 9827 2986 9840 3020
rect 8922 2957 8975 2972
rect 9783 2974 9840 2986
rect 9870 3186 9925 3198
rect 9870 3152 9883 3186
rect 9917 3174 9925 3186
rect 9991 3174 10044 3195
rect 9917 3152 9943 3174
rect 9870 3118 9943 3152
rect 9870 3084 9883 3118
rect 9917 3084 9943 3118
rect 9870 3050 9943 3084
rect 9870 3016 9883 3050
rect 9917 3016 9943 3050
rect 9870 2974 9943 3016
rect 9973 2995 10044 3174
rect 10074 3153 10127 3195
rect 10380 3182 10431 3194
rect 10380 3153 10388 3182
rect 10074 2995 10145 3153
rect 9973 2974 10026 2995
rect 10092 2953 10145 2995
rect 10175 3141 10235 3153
rect 10175 3107 10188 3141
rect 10222 3107 10235 3141
rect 10175 3073 10235 3107
rect 10175 3039 10188 3073
rect 10222 3039 10235 3073
rect 10175 3005 10235 3039
rect 10175 2971 10188 3005
rect 10222 2971 10235 3005
rect 10175 2953 10235 2971
rect 10265 3141 10332 3153
rect 10265 3107 10278 3141
rect 10312 3107 10332 3141
rect 10265 3049 10332 3107
rect 10265 3015 10278 3049
rect 10312 3015 10332 3049
rect 10265 2953 10332 3015
rect 10362 3148 10388 3153
rect 10422 3153 10431 3182
rect 11311 3186 11370 3198
rect 11000 3153 11119 3168
rect 10422 3148 10449 3153
rect 10362 2953 10449 3148
rect 10479 3114 10550 3153
rect 10479 3080 10492 3114
rect 10526 3080 10550 3114
rect 10479 2953 10550 3080
rect 10580 3117 10642 3153
rect 10580 3083 10593 3117
rect 10627 3083 10642 3117
rect 10580 2953 10642 3083
rect 10672 2953 10743 3153
rect 10773 3141 10833 3153
rect 10773 3107 10786 3141
rect 10820 3107 10833 3141
rect 10773 3030 10833 3107
rect 10773 2996 10786 3030
rect 10820 2996 10833 3030
rect 10773 2953 10833 2996
rect 10863 3141 10952 3153
rect 10863 3107 10905 3141
rect 10939 3107 10952 3141
rect 10863 3057 10952 3107
rect 10863 3023 10905 3057
rect 10939 3023 10952 3057
rect 10863 2953 10952 3023
rect 10982 3143 11119 3153
rect 10982 3109 10996 3143
rect 11030 3109 11071 3143
rect 11105 3109 11119 3143
rect 10982 2968 11119 3109
rect 11149 3156 11216 3168
rect 11149 3122 11170 3156
rect 11204 3122 11216 3156
rect 11149 3046 11216 3122
rect 11149 3012 11170 3046
rect 11204 3012 11216 3046
rect 11149 2968 11216 3012
rect 11311 3152 11323 3186
rect 11357 3152 11370 3186
rect 11311 3103 11370 3152
rect 11311 3069 11323 3103
rect 11357 3069 11370 3103
rect 11311 3020 11370 3069
rect 11311 2986 11323 3020
rect 11357 2986 11370 3020
rect 11311 2974 11370 2986
rect 11400 3186 11457 3198
rect 11400 3152 11413 3186
rect 11447 3152 11457 3186
rect 11400 3103 11457 3152
rect 11400 3069 11413 3103
rect 11447 3069 11457 3103
rect 11400 3020 11457 3069
rect 11400 2986 11413 3020
rect 11447 2986 11457 3020
rect 11400 2974 11457 2986
rect 11845 3182 11902 3194
rect 11845 3148 11855 3182
rect 11889 3148 11902 3182
rect 11845 3099 11902 3148
rect 11845 3065 11855 3099
rect 11889 3065 11902 3099
rect 11845 3016 11902 3065
rect 11845 2982 11855 3016
rect 11889 2982 11902 3016
rect 10982 2953 11035 2968
rect 11845 2970 11902 2982
rect 11932 3182 11987 3194
rect 11932 3148 11945 3182
rect 11979 3170 11987 3182
rect 12053 3170 12106 3191
rect 11979 3148 12005 3170
rect 11932 3114 12005 3148
rect 11932 3080 11945 3114
rect 11979 3080 12005 3114
rect 11932 3046 12005 3080
rect 11932 3012 11945 3046
rect 11979 3012 12005 3046
rect 11932 2970 12005 3012
rect 12035 2991 12106 3170
rect 12136 3149 12189 3191
rect 12442 3178 12493 3190
rect 12442 3149 12450 3178
rect 12136 2991 12207 3149
rect 12035 2970 12088 2991
rect 12154 2949 12207 2991
rect 12237 3137 12297 3149
rect 12237 3103 12250 3137
rect 12284 3103 12297 3137
rect 12237 3069 12297 3103
rect 12237 3035 12250 3069
rect 12284 3035 12297 3069
rect 12237 3001 12297 3035
rect 12237 2967 12250 3001
rect 12284 2967 12297 3001
rect 12237 2949 12297 2967
rect 12327 3137 12394 3149
rect 12327 3103 12340 3137
rect 12374 3103 12394 3137
rect 12327 3045 12394 3103
rect 12327 3011 12340 3045
rect 12374 3011 12394 3045
rect 12327 2949 12394 3011
rect 12424 3144 12450 3149
rect 12484 3149 12493 3178
rect 13373 3182 13432 3194
rect 13062 3149 13181 3164
rect 12484 3144 12511 3149
rect 12424 2949 12511 3144
rect 12541 3110 12612 3149
rect 12541 3076 12554 3110
rect 12588 3076 12612 3110
rect 12541 2949 12612 3076
rect 12642 3113 12704 3149
rect 12642 3079 12655 3113
rect 12689 3079 12704 3113
rect 12642 2949 12704 3079
rect 12734 2949 12805 3149
rect 12835 3137 12895 3149
rect 12835 3103 12848 3137
rect 12882 3103 12895 3137
rect 12835 3026 12895 3103
rect 12835 2992 12848 3026
rect 12882 2992 12895 3026
rect 12835 2949 12895 2992
rect 12925 3137 13014 3149
rect 12925 3103 12967 3137
rect 13001 3103 13014 3137
rect 12925 3053 13014 3103
rect 12925 3019 12967 3053
rect 13001 3019 13014 3053
rect 12925 2949 13014 3019
rect 13044 3139 13181 3149
rect 13044 3105 13058 3139
rect 13092 3105 13133 3139
rect 13167 3105 13181 3139
rect 13044 2964 13181 3105
rect 13211 3152 13278 3164
rect 13211 3118 13232 3152
rect 13266 3118 13278 3152
rect 13211 3042 13278 3118
rect 13211 3008 13232 3042
rect 13266 3008 13278 3042
rect 13211 2964 13278 3008
rect 13373 3148 13385 3182
rect 13419 3148 13432 3182
rect 13373 3099 13432 3148
rect 13373 3065 13385 3099
rect 13419 3065 13432 3099
rect 13373 3016 13432 3065
rect 13373 2982 13385 3016
rect 13419 2982 13432 3016
rect 13373 2970 13432 2982
rect 13462 3182 13519 3194
rect 13462 3148 13475 3182
rect 13509 3148 13519 3182
rect 13462 3099 13519 3148
rect 13462 3065 13475 3099
rect 13509 3065 13519 3099
rect 13462 3016 13519 3065
rect 13462 2982 13475 3016
rect 13509 2982 13519 3016
rect 13462 2970 13519 2982
rect 13919 3180 13976 3192
rect 13919 3146 13929 3180
rect 13963 3146 13976 3180
rect 13919 3097 13976 3146
rect 13919 3063 13929 3097
rect 13963 3063 13976 3097
rect 13919 3014 13976 3063
rect 13919 2980 13929 3014
rect 13963 2980 13976 3014
rect 13044 2949 13097 2964
rect 13919 2968 13976 2980
rect 14006 3180 14061 3192
rect 14006 3146 14019 3180
rect 14053 3168 14061 3180
rect 14127 3168 14180 3189
rect 14053 3146 14079 3168
rect 14006 3112 14079 3146
rect 14006 3078 14019 3112
rect 14053 3078 14079 3112
rect 14006 3044 14079 3078
rect 14006 3010 14019 3044
rect 14053 3010 14079 3044
rect 14006 2968 14079 3010
rect 14109 2989 14180 3168
rect 14210 3147 14263 3189
rect 14516 3176 14567 3188
rect 14516 3147 14524 3176
rect 14210 2989 14281 3147
rect 14109 2968 14162 2989
rect 14228 2947 14281 2989
rect 14311 3135 14371 3147
rect 14311 3101 14324 3135
rect 14358 3101 14371 3135
rect 14311 3067 14371 3101
rect 14311 3033 14324 3067
rect 14358 3033 14371 3067
rect 14311 2999 14371 3033
rect 14311 2965 14324 2999
rect 14358 2965 14371 2999
rect 14311 2947 14371 2965
rect 14401 3135 14468 3147
rect 14401 3101 14414 3135
rect 14448 3101 14468 3135
rect 14401 3043 14468 3101
rect 14401 3009 14414 3043
rect 14448 3009 14468 3043
rect 14401 2947 14468 3009
rect 14498 3142 14524 3147
rect 14558 3147 14567 3176
rect 15447 3180 15506 3192
rect 15136 3147 15255 3162
rect 14558 3142 14585 3147
rect 14498 2947 14585 3142
rect 14615 3108 14686 3147
rect 14615 3074 14628 3108
rect 14662 3074 14686 3108
rect 14615 2947 14686 3074
rect 14716 3111 14778 3147
rect 14716 3077 14729 3111
rect 14763 3077 14778 3111
rect 14716 2947 14778 3077
rect 14808 2947 14879 3147
rect 14909 3135 14969 3147
rect 14909 3101 14922 3135
rect 14956 3101 14969 3135
rect 14909 3024 14969 3101
rect 14909 2990 14922 3024
rect 14956 2990 14969 3024
rect 14909 2947 14969 2990
rect 14999 3135 15088 3147
rect 14999 3101 15041 3135
rect 15075 3101 15088 3135
rect 14999 3051 15088 3101
rect 14999 3017 15041 3051
rect 15075 3017 15088 3051
rect 14999 2947 15088 3017
rect 15118 3137 15255 3147
rect 15118 3103 15132 3137
rect 15166 3103 15207 3137
rect 15241 3103 15255 3137
rect 15118 2962 15255 3103
rect 15285 3150 15352 3162
rect 15285 3116 15306 3150
rect 15340 3116 15352 3150
rect 15285 3040 15352 3116
rect 15285 3006 15306 3040
rect 15340 3006 15352 3040
rect 15285 2962 15352 3006
rect 15447 3146 15459 3180
rect 15493 3146 15506 3180
rect 15447 3097 15506 3146
rect 15447 3063 15459 3097
rect 15493 3063 15506 3097
rect 15447 3014 15506 3063
rect 15447 2980 15459 3014
rect 15493 2980 15506 3014
rect 15447 2968 15506 2980
rect 15536 3180 15593 3192
rect 15536 3146 15549 3180
rect 15583 3146 15593 3180
rect 15536 3097 15593 3146
rect 15536 3063 15549 3097
rect 15583 3063 15593 3097
rect 15536 3014 15593 3063
rect 15536 2980 15549 3014
rect 15583 2980 15593 3014
rect 15536 2968 15593 2980
rect 15981 3176 16038 3188
rect 15981 3142 15991 3176
rect 16025 3142 16038 3176
rect 15981 3093 16038 3142
rect 15981 3059 15991 3093
rect 16025 3059 16038 3093
rect 15981 3010 16038 3059
rect 15981 2976 15991 3010
rect 16025 2976 16038 3010
rect 15118 2947 15171 2962
rect 15981 2964 16038 2976
rect 16068 3176 16123 3188
rect 16068 3142 16081 3176
rect 16115 3164 16123 3176
rect 16189 3164 16242 3185
rect 16115 3142 16141 3164
rect 16068 3108 16141 3142
rect 16068 3074 16081 3108
rect 16115 3074 16141 3108
rect 16068 3040 16141 3074
rect 16068 3006 16081 3040
rect 16115 3006 16141 3040
rect 16068 2964 16141 3006
rect 16171 2985 16242 3164
rect 16272 3143 16325 3185
rect 16578 3172 16629 3184
rect 16578 3143 16586 3172
rect 16272 2985 16343 3143
rect 16171 2964 16224 2985
rect 16290 2943 16343 2985
rect 16373 3131 16433 3143
rect 16373 3097 16386 3131
rect 16420 3097 16433 3131
rect 16373 3063 16433 3097
rect 16373 3029 16386 3063
rect 16420 3029 16433 3063
rect 16373 2995 16433 3029
rect 16373 2961 16386 2995
rect 16420 2961 16433 2995
rect 16373 2943 16433 2961
rect 16463 3131 16530 3143
rect 16463 3097 16476 3131
rect 16510 3097 16530 3131
rect 16463 3039 16530 3097
rect 16463 3005 16476 3039
rect 16510 3005 16530 3039
rect 16463 2943 16530 3005
rect 16560 3138 16586 3143
rect 16620 3143 16629 3172
rect 17509 3176 17568 3188
rect 17198 3143 17317 3158
rect 16620 3138 16647 3143
rect 16560 2943 16647 3138
rect 16677 3104 16748 3143
rect 16677 3070 16690 3104
rect 16724 3070 16748 3104
rect 16677 2943 16748 3070
rect 16778 3107 16840 3143
rect 16778 3073 16791 3107
rect 16825 3073 16840 3107
rect 16778 2943 16840 3073
rect 16870 2943 16941 3143
rect 16971 3131 17031 3143
rect 16971 3097 16984 3131
rect 17018 3097 17031 3131
rect 16971 3020 17031 3097
rect 16971 2986 16984 3020
rect 17018 2986 17031 3020
rect 16971 2943 17031 2986
rect 17061 3131 17150 3143
rect 17061 3097 17103 3131
rect 17137 3097 17150 3131
rect 17061 3047 17150 3097
rect 17061 3013 17103 3047
rect 17137 3013 17150 3047
rect 17061 2943 17150 3013
rect 17180 3133 17317 3143
rect 17180 3099 17194 3133
rect 17228 3099 17269 3133
rect 17303 3099 17317 3133
rect 17180 2958 17317 3099
rect 17347 3146 17414 3158
rect 17347 3112 17368 3146
rect 17402 3112 17414 3146
rect 17347 3036 17414 3112
rect 17347 3002 17368 3036
rect 17402 3002 17414 3036
rect 17347 2958 17414 3002
rect 17509 3142 17521 3176
rect 17555 3142 17568 3176
rect 17509 3093 17568 3142
rect 17509 3059 17521 3093
rect 17555 3059 17568 3093
rect 17509 3010 17568 3059
rect 17509 2976 17521 3010
rect 17555 2976 17568 3010
rect 17509 2964 17568 2976
rect 17598 3176 17655 3188
rect 17598 3142 17611 3176
rect 17645 3142 17655 3176
rect 17598 3093 17655 3142
rect 17598 3059 17611 3093
rect 17645 3059 17655 3093
rect 17598 3010 17655 3059
rect 17598 2976 17611 3010
rect 17645 2976 17655 3010
rect 17598 2964 17655 2976
rect 22612 3071 22664 3083
rect 22612 3037 22620 3071
rect 22654 3037 22664 3071
rect 22612 3003 22664 3037
rect 22612 2969 22620 3003
rect 22654 2969 22664 3003
rect 17180 2943 17233 2958
rect 22612 2935 22664 2969
rect 22612 2901 22620 2935
rect 22654 2901 22664 2935
rect 22612 2883 22664 2901
rect 22694 3071 22746 3083
rect 22694 3037 22704 3071
rect 22738 3037 22746 3071
rect 22694 3003 22746 3037
rect 22694 2969 22704 3003
rect 22738 2969 22746 3003
rect 22694 2935 22746 2969
rect 22694 2901 22704 2935
rect 22738 2901 22746 2935
rect 22694 2883 22746 2901
rect 23197 3069 23249 3081
rect 23197 3035 23205 3069
rect 23239 3035 23249 3069
rect 23197 3001 23249 3035
rect 23197 2967 23205 3001
rect 23239 2967 23249 3001
rect 23197 2933 23249 2967
rect 23197 2899 23205 2933
rect 23239 2899 23249 2933
rect 23197 2881 23249 2899
rect 23279 3069 23333 3081
rect 23279 3035 23289 3069
rect 23323 3035 23333 3069
rect 23279 3001 23333 3035
rect 23279 2967 23289 3001
rect 23323 2967 23333 3001
rect 23279 2933 23333 2967
rect 23279 2899 23289 2933
rect 23323 2899 23333 2933
rect 23279 2881 23333 2899
rect 23363 3069 23415 3081
rect 23363 3035 23373 3069
rect 23407 3035 23415 3069
rect 23363 3001 23415 3035
rect 23363 2967 23373 3001
rect 23407 2967 23415 3001
rect 23363 2933 23415 2967
rect 23363 2899 23373 2933
rect 23407 2899 23415 2933
rect 23363 2881 23415 2899
rect 23813 3057 23865 3069
rect 23813 3023 23821 3057
rect 23855 3023 23865 3057
rect 23813 2989 23865 3023
rect 23813 2955 23821 2989
rect 23855 2955 23865 2989
rect 23813 2921 23865 2955
rect 23813 2887 23821 2921
rect 23855 2887 23865 2921
rect 23813 2869 23865 2887
rect 23895 3057 23949 3069
rect 23895 3023 23905 3057
rect 23939 3023 23949 3057
rect 23895 2989 23949 3023
rect 23895 2955 23905 2989
rect 23939 2955 23949 2989
rect 23895 2921 23949 2955
rect 23895 2887 23905 2921
rect 23939 2887 23949 2921
rect 23895 2869 23949 2887
rect 23979 3057 24033 3069
rect 23979 3023 23989 3057
rect 24023 3023 24033 3057
rect 23979 2989 24033 3023
rect 23979 2955 23989 2989
rect 24023 2955 24033 2989
rect 23979 2869 24033 2955
rect 24063 3057 24117 3069
rect 24063 3023 24073 3057
rect 24107 3023 24117 3057
rect 24063 2989 24117 3023
rect 24063 2955 24073 2989
rect 24107 2955 24117 2989
rect 24063 2921 24117 2955
rect 24063 2887 24073 2921
rect 24107 2887 24117 2921
rect 24063 2869 24117 2887
rect 24147 3057 24199 3069
rect 24147 3023 24157 3057
rect 24191 3023 24199 3057
rect 24147 2869 24199 3023
rect 24627 3043 24713 3055
rect 24627 3009 24635 3043
rect 24669 3009 24713 3043
rect 24627 2975 24713 3009
rect 24627 2941 24635 2975
rect 24669 2941 24713 2975
rect 24627 2907 24713 2941
rect 24627 2873 24635 2907
rect 24669 2873 24713 2907
rect 24627 2855 24713 2873
rect 24743 3043 24797 3055
rect 24743 3009 24753 3043
rect 24787 3009 24797 3043
rect 24743 2975 24797 3009
rect 24743 2941 24753 2975
rect 24787 2941 24797 2975
rect 24743 2907 24797 2941
rect 24743 2873 24753 2907
rect 24787 2873 24797 2907
rect 24743 2855 24797 2873
rect 24827 3043 24881 3055
rect 24827 3009 24837 3043
rect 24871 3009 24881 3043
rect 24827 2975 24881 3009
rect 24827 2941 24837 2975
rect 24871 2941 24881 2975
rect 24827 2855 24881 2941
rect 24911 3043 24965 3055
rect 24911 3009 24921 3043
rect 24955 3009 24965 3043
rect 24911 2975 24965 3009
rect 24911 2941 24921 2975
rect 24955 2941 24965 2975
rect 24911 2907 24965 2941
rect 24911 2873 24921 2907
rect 24955 2873 24965 2907
rect 24911 2855 24965 2873
rect 24995 3043 25049 3055
rect 24995 3009 25005 3043
rect 25039 3009 25049 3043
rect 24995 2975 25049 3009
rect 24995 2941 25005 2975
rect 25039 2941 25049 2975
rect 24995 2855 25049 2941
rect 25079 3043 25133 3055
rect 25079 3009 25089 3043
rect 25123 3009 25133 3043
rect 25079 2975 25133 3009
rect 25079 2941 25089 2975
rect 25123 2941 25133 2975
rect 25079 2907 25133 2941
rect 25079 2873 25089 2907
rect 25123 2873 25133 2907
rect 25079 2855 25133 2873
rect 25163 3043 25217 3055
rect 25163 3009 25173 3043
rect 25207 3009 25217 3043
rect 25163 2855 25217 3009
<< ndiffc >>
rect 8138 4332 8172 4366
rect 8138 4242 8172 4276
rect 8224 4332 8258 4366
rect 8224 4242 8258 4276
rect 8310 4332 8344 4366
rect 8310 4242 8344 4276
rect 1537 2796 1571 2830
rect 1537 2706 1571 2740
rect 1641 2668 1675 2702
rect 1902 2713 1936 2747
rect 2018 2720 2052 2754
rect 2128 2668 2162 2702
rect 2230 2720 2264 2754
rect 2344 2712 2378 2746
rect 2523 2723 2557 2757
rect 2625 2671 2659 2705
rect 2719 2671 2753 2705
rect 2864 2664 2898 2698
rect 2966 2732 3000 2766
rect 3070 2724 3104 2758
rect 3156 2796 3190 2830
rect 3156 2706 3190 2740
rect 3599 2792 3633 2826
rect 3599 2702 3633 2736
rect 3703 2664 3737 2698
rect 3964 2709 3998 2743
rect 4080 2716 4114 2750
rect 4190 2664 4224 2698
rect 4292 2716 4326 2750
rect 4406 2708 4440 2742
rect 4585 2719 4619 2753
rect 4687 2667 4721 2701
rect 4781 2667 4815 2701
rect 4926 2660 4960 2694
rect 5028 2728 5062 2762
rect 5132 2720 5166 2754
rect 5218 2792 5252 2826
rect 5218 2702 5252 2736
rect 5673 2790 5707 2824
rect 5673 2700 5707 2734
rect 5777 2662 5811 2696
rect 6038 2707 6072 2741
rect 6154 2714 6188 2748
rect 6264 2662 6298 2696
rect 6366 2714 6400 2748
rect 6480 2706 6514 2740
rect 6659 2717 6693 2751
rect 6761 2665 6795 2699
rect 6855 2665 6889 2699
rect 7000 2658 7034 2692
rect 7102 2726 7136 2760
rect 7206 2718 7240 2752
rect 7292 2790 7326 2824
rect 7292 2700 7326 2734
rect 7735 2786 7769 2820
rect 7735 2696 7769 2730
rect 7839 2658 7873 2692
rect 8100 2703 8134 2737
rect 8216 2710 8250 2744
rect 8326 2658 8360 2692
rect 8428 2710 8462 2744
rect 8542 2702 8576 2736
rect 8721 2713 8755 2747
rect 8823 2661 8857 2695
rect 8917 2661 8951 2695
rect 9062 2654 9096 2688
rect 9164 2722 9198 2756
rect 9268 2714 9302 2748
rect 9354 2786 9388 2820
rect 9354 2696 9388 2730
rect 9795 2782 9829 2816
rect 9795 2692 9829 2726
rect 9899 2654 9933 2688
rect 10160 2699 10194 2733
rect 10276 2706 10310 2740
rect 10386 2654 10420 2688
rect 10488 2706 10522 2740
rect 10602 2698 10636 2732
rect 10781 2709 10815 2743
rect 10883 2657 10917 2691
rect 10977 2657 11011 2691
rect 11122 2650 11156 2684
rect 11224 2718 11258 2752
rect 11328 2710 11362 2744
rect 11414 2782 11448 2816
rect 11414 2692 11448 2726
rect 11857 2778 11891 2812
rect 11857 2688 11891 2722
rect 11961 2650 11995 2684
rect 12222 2695 12256 2729
rect 12338 2702 12372 2736
rect 12448 2650 12482 2684
rect 12550 2702 12584 2736
rect 12664 2694 12698 2728
rect 12843 2705 12877 2739
rect 12945 2653 12979 2687
rect 13039 2653 13073 2687
rect 13184 2646 13218 2680
rect 13286 2714 13320 2748
rect 13390 2706 13424 2740
rect 13476 2778 13510 2812
rect 13476 2688 13510 2722
rect 13931 2776 13965 2810
rect 13931 2686 13965 2720
rect 14035 2648 14069 2682
rect 14296 2693 14330 2727
rect 14412 2700 14446 2734
rect 14522 2648 14556 2682
rect 14624 2700 14658 2734
rect 14738 2692 14772 2726
rect 14917 2703 14951 2737
rect 15019 2651 15053 2685
rect 15113 2651 15147 2685
rect 15258 2644 15292 2678
rect 15360 2712 15394 2746
rect 15464 2704 15498 2738
rect 15550 2776 15584 2810
rect 15550 2686 15584 2720
rect 15993 2772 16027 2806
rect 15993 2682 16027 2716
rect 16097 2644 16131 2678
rect 16358 2689 16392 2723
rect 16474 2696 16508 2730
rect 16584 2644 16618 2678
rect 16686 2696 16720 2730
rect 16800 2688 16834 2722
rect 16979 2699 17013 2733
rect 17081 2647 17115 2681
rect 17175 2647 17209 2681
rect 17320 2640 17354 2674
rect 17422 2708 17456 2742
rect 17526 2700 17560 2734
rect 17612 2772 17646 2806
rect 17612 2682 17646 2716
rect 22620 2717 22654 2751
rect 22620 2649 22654 2683
rect 22704 2717 22738 2751
rect 22704 2649 22738 2683
rect 23205 2715 23239 2749
rect 23205 2643 23239 2677
rect 23289 2715 23323 2749
rect 23289 2643 23323 2677
rect 23373 2715 23407 2749
rect 23373 2643 23407 2677
rect 23821 2631 23855 2665
rect 23905 2639 23939 2673
rect 23989 2631 24023 2665
rect 24073 2639 24107 2673
rect 24157 2632 24191 2666
rect 24645 2617 24679 2651
rect 24753 2625 24787 2659
rect 24837 2617 24871 2651
rect 24921 2625 24955 2659
rect 25005 2617 25039 2651
rect 25089 2625 25123 2659
rect 25173 2618 25207 2652
<< pdiffc >>
rect 8135 4038 8169 4072
rect 8135 3955 8169 3989
rect 8135 3872 8169 3906
rect 8225 4038 8259 4072
rect 8225 3955 8259 3989
rect 8225 3872 8259 3906
rect 8315 4012 8349 4046
rect 8315 3942 8349 3976
rect 8315 3872 8349 3906
rect 1535 3166 1569 3200
rect 1535 3083 1569 3117
rect 1535 3000 1569 3034
rect 1625 3166 1659 3200
rect 1625 3098 1659 3132
rect 1625 3030 1659 3064
rect 1930 3121 1964 3155
rect 1930 3053 1964 3087
rect 1930 2985 1964 3019
rect 2020 3121 2054 3155
rect 2020 3029 2054 3063
rect 2130 3162 2164 3196
rect 2234 3094 2268 3128
rect 2335 3097 2369 3131
rect 2528 3121 2562 3155
rect 2528 3010 2562 3044
rect 2647 3121 2681 3155
rect 2647 3037 2681 3071
rect 2738 3123 2772 3157
rect 2813 3123 2847 3157
rect 2912 3136 2946 3170
rect 2912 3026 2946 3060
rect 3065 3166 3099 3200
rect 3065 3083 3099 3117
rect 3065 3000 3099 3034
rect 3155 3166 3189 3200
rect 3155 3083 3189 3117
rect 3155 3000 3189 3034
rect 3597 3162 3631 3196
rect 3597 3079 3631 3113
rect 3597 2996 3631 3030
rect 3687 3162 3721 3196
rect 3687 3094 3721 3128
rect 3687 3026 3721 3060
rect 3992 3117 4026 3151
rect 3992 3049 4026 3083
rect 3992 2981 4026 3015
rect 4082 3117 4116 3151
rect 4082 3025 4116 3059
rect 4192 3158 4226 3192
rect 4296 3090 4330 3124
rect 4397 3093 4431 3127
rect 4590 3117 4624 3151
rect 4590 3006 4624 3040
rect 4709 3117 4743 3151
rect 4709 3033 4743 3067
rect 4800 3119 4834 3153
rect 4875 3119 4909 3153
rect 4974 3132 5008 3166
rect 4974 3022 5008 3056
rect 5127 3162 5161 3196
rect 5127 3079 5161 3113
rect 5127 2996 5161 3030
rect 5217 3162 5251 3196
rect 5217 3079 5251 3113
rect 5217 2996 5251 3030
rect 5671 3160 5705 3194
rect 5671 3077 5705 3111
rect 5671 2994 5705 3028
rect 5761 3160 5795 3194
rect 5761 3092 5795 3126
rect 5761 3024 5795 3058
rect 6066 3115 6100 3149
rect 6066 3047 6100 3081
rect 6066 2979 6100 3013
rect 6156 3115 6190 3149
rect 6156 3023 6190 3057
rect 6266 3156 6300 3190
rect 6370 3088 6404 3122
rect 6471 3091 6505 3125
rect 6664 3115 6698 3149
rect 6664 3004 6698 3038
rect 6783 3115 6817 3149
rect 6783 3031 6817 3065
rect 6874 3117 6908 3151
rect 6949 3117 6983 3151
rect 7048 3130 7082 3164
rect 7048 3020 7082 3054
rect 7201 3160 7235 3194
rect 7201 3077 7235 3111
rect 7201 2994 7235 3028
rect 7291 3160 7325 3194
rect 7291 3077 7325 3111
rect 7291 2994 7325 3028
rect 7733 3156 7767 3190
rect 7733 3073 7767 3107
rect 7733 2990 7767 3024
rect 7823 3156 7857 3190
rect 7823 3088 7857 3122
rect 7823 3020 7857 3054
rect 8128 3111 8162 3145
rect 8128 3043 8162 3077
rect 8128 2975 8162 3009
rect 8218 3111 8252 3145
rect 8218 3019 8252 3053
rect 8328 3152 8362 3186
rect 8432 3084 8466 3118
rect 8533 3087 8567 3121
rect 8726 3111 8760 3145
rect 8726 3000 8760 3034
rect 8845 3111 8879 3145
rect 8845 3027 8879 3061
rect 8936 3113 8970 3147
rect 9011 3113 9045 3147
rect 9110 3126 9144 3160
rect 9110 3016 9144 3050
rect 9263 3156 9297 3190
rect 9263 3073 9297 3107
rect 9263 2990 9297 3024
rect 9353 3156 9387 3190
rect 9353 3073 9387 3107
rect 9353 2990 9387 3024
rect 9793 3152 9827 3186
rect 9793 3069 9827 3103
rect 9793 2986 9827 3020
rect 9883 3152 9917 3186
rect 9883 3084 9917 3118
rect 9883 3016 9917 3050
rect 10188 3107 10222 3141
rect 10188 3039 10222 3073
rect 10188 2971 10222 3005
rect 10278 3107 10312 3141
rect 10278 3015 10312 3049
rect 10388 3148 10422 3182
rect 10492 3080 10526 3114
rect 10593 3083 10627 3117
rect 10786 3107 10820 3141
rect 10786 2996 10820 3030
rect 10905 3107 10939 3141
rect 10905 3023 10939 3057
rect 10996 3109 11030 3143
rect 11071 3109 11105 3143
rect 11170 3122 11204 3156
rect 11170 3012 11204 3046
rect 11323 3152 11357 3186
rect 11323 3069 11357 3103
rect 11323 2986 11357 3020
rect 11413 3152 11447 3186
rect 11413 3069 11447 3103
rect 11413 2986 11447 3020
rect 11855 3148 11889 3182
rect 11855 3065 11889 3099
rect 11855 2982 11889 3016
rect 11945 3148 11979 3182
rect 11945 3080 11979 3114
rect 11945 3012 11979 3046
rect 12250 3103 12284 3137
rect 12250 3035 12284 3069
rect 12250 2967 12284 3001
rect 12340 3103 12374 3137
rect 12340 3011 12374 3045
rect 12450 3144 12484 3178
rect 12554 3076 12588 3110
rect 12655 3079 12689 3113
rect 12848 3103 12882 3137
rect 12848 2992 12882 3026
rect 12967 3103 13001 3137
rect 12967 3019 13001 3053
rect 13058 3105 13092 3139
rect 13133 3105 13167 3139
rect 13232 3118 13266 3152
rect 13232 3008 13266 3042
rect 13385 3148 13419 3182
rect 13385 3065 13419 3099
rect 13385 2982 13419 3016
rect 13475 3148 13509 3182
rect 13475 3065 13509 3099
rect 13475 2982 13509 3016
rect 13929 3146 13963 3180
rect 13929 3063 13963 3097
rect 13929 2980 13963 3014
rect 14019 3146 14053 3180
rect 14019 3078 14053 3112
rect 14019 3010 14053 3044
rect 14324 3101 14358 3135
rect 14324 3033 14358 3067
rect 14324 2965 14358 2999
rect 14414 3101 14448 3135
rect 14414 3009 14448 3043
rect 14524 3142 14558 3176
rect 14628 3074 14662 3108
rect 14729 3077 14763 3111
rect 14922 3101 14956 3135
rect 14922 2990 14956 3024
rect 15041 3101 15075 3135
rect 15041 3017 15075 3051
rect 15132 3103 15166 3137
rect 15207 3103 15241 3137
rect 15306 3116 15340 3150
rect 15306 3006 15340 3040
rect 15459 3146 15493 3180
rect 15459 3063 15493 3097
rect 15459 2980 15493 3014
rect 15549 3146 15583 3180
rect 15549 3063 15583 3097
rect 15549 2980 15583 3014
rect 15991 3142 16025 3176
rect 15991 3059 16025 3093
rect 15991 2976 16025 3010
rect 16081 3142 16115 3176
rect 16081 3074 16115 3108
rect 16081 3006 16115 3040
rect 16386 3097 16420 3131
rect 16386 3029 16420 3063
rect 16386 2961 16420 2995
rect 16476 3097 16510 3131
rect 16476 3005 16510 3039
rect 16586 3138 16620 3172
rect 16690 3070 16724 3104
rect 16791 3073 16825 3107
rect 16984 3097 17018 3131
rect 16984 2986 17018 3020
rect 17103 3097 17137 3131
rect 17103 3013 17137 3047
rect 17194 3099 17228 3133
rect 17269 3099 17303 3133
rect 17368 3112 17402 3146
rect 17368 3002 17402 3036
rect 17521 3142 17555 3176
rect 17521 3059 17555 3093
rect 17521 2976 17555 3010
rect 17611 3142 17645 3176
rect 17611 3059 17645 3093
rect 17611 2976 17645 3010
rect 22620 3037 22654 3071
rect 22620 2969 22654 3003
rect 22620 2901 22654 2935
rect 22704 3037 22738 3071
rect 22704 2969 22738 3003
rect 22704 2901 22738 2935
rect 23205 3035 23239 3069
rect 23205 2967 23239 3001
rect 23205 2899 23239 2933
rect 23289 3035 23323 3069
rect 23289 2967 23323 3001
rect 23289 2899 23323 2933
rect 23373 3035 23407 3069
rect 23373 2967 23407 3001
rect 23373 2899 23407 2933
rect 23821 3023 23855 3057
rect 23821 2955 23855 2989
rect 23821 2887 23855 2921
rect 23905 3023 23939 3057
rect 23905 2955 23939 2989
rect 23905 2887 23939 2921
rect 23989 3023 24023 3057
rect 23989 2955 24023 2989
rect 24073 3023 24107 3057
rect 24073 2955 24107 2989
rect 24073 2887 24107 2921
rect 24157 3023 24191 3057
rect 24635 3009 24669 3043
rect 24635 2941 24669 2975
rect 24635 2873 24669 2907
rect 24753 3009 24787 3043
rect 24753 2941 24787 2975
rect 24753 2873 24787 2907
rect 24837 3009 24871 3043
rect 24837 2941 24871 2975
rect 24921 3009 24955 3043
rect 24921 2941 24955 2975
rect 24921 2873 24955 2907
rect 25005 3009 25039 3043
rect 25005 2941 25039 2975
rect 25089 3009 25123 3043
rect 25089 2941 25123 2975
rect 25089 2873 25123 2907
rect 25173 3009 25207 3043
<< poly >>
rect 8183 4378 8213 4404
rect 8269 4378 8299 4404
rect 8183 4192 8213 4230
rect 8269 4192 8299 4230
rect 8179 4176 8365 4192
rect 8179 4162 8315 4176
rect 8179 4099 8215 4162
rect 8269 4142 8315 4162
rect 8349 4142 8365 4176
rect 8269 4126 8365 4142
rect 8269 4099 8305 4126
rect 8182 4084 8212 4099
rect 8272 4084 8302 4099
rect 8182 3834 8212 3860
rect 8272 3834 8302 3860
rect 1582 3212 1612 3238
rect 1783 3235 2894 3265
rect 1783 3224 1819 3235
rect 1685 3188 1715 3214
rect 1786 3209 1816 3224
rect 1887 3167 1917 3193
rect 1977 3167 2007 3193
rect 2071 3182 2107 3235
rect 2074 3167 2104 3182
rect 1786 2994 1816 3009
rect 1582 2973 1612 2988
rect 1685 2973 1715 2988
rect 1579 2946 1615 2973
rect 1567 2930 1633 2946
rect 1682 2930 1718 2973
rect 1783 2963 1819 2994
rect 2191 3167 2221 3193
rect 2292 3167 2322 3193
rect 2384 3167 2414 3193
rect 2482 3182 2518 3235
rect 2858 3197 2894 3235
rect 3112 3212 3142 3238
rect 2485 3167 2515 3182
rect 2575 3167 2605 3193
rect 2694 3167 2724 3193
rect 2861 3182 2891 3197
rect 3644 3208 3674 3234
rect 3845 3231 4956 3261
rect 3845 3220 3881 3231
rect 2861 2967 2891 2982
rect 3112 2973 3142 2988
rect 3747 3184 3777 3210
rect 3848 3205 3878 3220
rect 3949 3163 3979 3189
rect 4039 3163 4069 3189
rect 4133 3178 4169 3231
rect 4136 3163 4166 3178
rect 3848 2990 3878 3005
rect 1567 2896 1583 2930
rect 1617 2896 1633 2930
rect 1567 2880 1633 2896
rect 1675 2914 1741 2930
rect 1675 2880 1691 2914
rect 1725 2880 1741 2914
rect 1582 2842 1612 2880
rect 1675 2864 1741 2880
rect 1705 2823 1735 2864
rect 1783 2823 1813 2963
rect 1887 2952 1917 2967
rect 1977 2952 2007 2967
rect 2074 2952 2104 2967
rect 2191 2952 2221 2967
rect 2292 2952 2322 2967
rect 2384 2952 2414 2967
rect 2485 2952 2515 2967
rect 2575 2952 2605 2967
rect 2694 2952 2724 2967
rect 1884 2935 1920 2952
rect 1974 2935 2010 2952
rect 1855 2919 1921 2935
rect 1855 2885 1871 2919
rect 1905 2885 1921 2919
rect 1855 2869 1921 2885
rect 1963 2919 2029 2935
rect 1963 2885 1979 2919
rect 2013 2885 2029 2919
rect 1963 2869 2029 2885
rect 1861 2823 1891 2869
rect 1969 2823 1999 2869
rect 2071 2838 2107 2952
rect 2188 2911 2224 2952
rect 2289 2935 2325 2952
rect 2158 2895 2224 2911
rect 2158 2861 2174 2895
rect 2208 2861 2224 2895
rect 2266 2919 2332 2935
rect 2266 2885 2282 2919
rect 2316 2885 2332 2919
rect 2381 2911 2417 2952
rect 2266 2869 2332 2885
rect 2374 2895 2440 2911
rect 2158 2845 2224 2861
rect 2071 2823 2101 2838
rect 2189 2823 2219 2845
rect 2275 2823 2305 2869
rect 2374 2861 2390 2895
rect 2424 2861 2440 2895
rect 2374 2845 2440 2861
rect 2404 2823 2434 2845
rect 2482 2838 2518 2952
rect 2572 2935 2608 2952
rect 2691 2935 2727 2952
rect 2858 2950 2894 2967
rect 2560 2919 2626 2935
rect 2560 2885 2576 2919
rect 2610 2885 2626 2919
rect 2560 2869 2626 2885
rect 2674 2919 2740 2935
rect 2674 2885 2690 2919
rect 2724 2885 2740 2919
rect 2674 2872 2740 2885
rect 2858 2934 2992 2950
rect 2858 2900 2874 2934
rect 2908 2900 2942 2934
rect 2976 2900 2992 2934
rect 3109 2930 3145 2973
rect 3644 2969 3674 2984
rect 3747 2969 3777 2984
rect 3641 2942 3677 2969
rect 2858 2884 2992 2900
rect 3040 2914 3145 2930
rect 2482 2823 2512 2838
rect 2568 2823 2598 2869
rect 2674 2842 2810 2872
rect 2780 2823 2810 2842
rect 2925 2823 2955 2884
rect 3040 2880 3056 2914
rect 3090 2880 3145 2914
rect 3040 2864 3145 2880
rect 3629 2926 3695 2942
rect 3744 2926 3780 2969
rect 3845 2959 3881 2990
rect 4253 3163 4283 3189
rect 4354 3163 4384 3189
rect 4446 3163 4476 3189
rect 4544 3178 4580 3231
rect 4920 3193 4956 3231
rect 5174 3208 5204 3234
rect 4547 3163 4577 3178
rect 4637 3163 4667 3189
rect 4756 3163 4786 3189
rect 4923 3178 4953 3193
rect 5718 3206 5748 3232
rect 5919 3229 7030 3259
rect 5919 3218 5955 3229
rect 4923 2963 4953 2978
rect 5174 2969 5204 2984
rect 5821 3182 5851 3208
rect 5922 3203 5952 3218
rect 6023 3161 6053 3187
rect 6113 3161 6143 3187
rect 6207 3176 6243 3229
rect 6210 3161 6240 3176
rect 5922 2988 5952 3003
rect 3629 2892 3645 2926
rect 3679 2892 3695 2926
rect 3629 2876 3695 2892
rect 3737 2910 3803 2926
rect 3737 2876 3753 2910
rect 3787 2876 3803 2910
rect 3115 2842 3145 2864
rect 1582 2668 1612 2694
rect 1705 2669 1735 2695
rect 1783 2669 1813 2695
rect 1861 2669 1891 2695
rect 1969 2669 1999 2695
rect 2071 2669 2101 2695
rect 2189 2669 2219 2695
rect 2275 2669 2305 2695
rect 2404 2669 2434 2695
rect 2482 2669 2512 2695
rect 2568 2669 2598 2695
rect 2780 2669 2810 2695
rect 2925 2669 2955 2695
rect 3644 2838 3674 2876
rect 3737 2860 3803 2876
rect 3115 2668 3145 2694
rect 3767 2819 3797 2860
rect 3845 2819 3875 2959
rect 3949 2948 3979 2963
rect 4039 2948 4069 2963
rect 4136 2948 4166 2963
rect 4253 2948 4283 2963
rect 4354 2948 4384 2963
rect 4446 2948 4476 2963
rect 4547 2948 4577 2963
rect 4637 2948 4667 2963
rect 4756 2948 4786 2963
rect 3946 2931 3982 2948
rect 4036 2931 4072 2948
rect 3917 2915 3983 2931
rect 3917 2881 3933 2915
rect 3967 2881 3983 2915
rect 3917 2865 3983 2881
rect 4025 2915 4091 2931
rect 4025 2881 4041 2915
rect 4075 2881 4091 2915
rect 4025 2865 4091 2881
rect 3923 2819 3953 2865
rect 4031 2819 4061 2865
rect 4133 2834 4169 2948
rect 4250 2907 4286 2948
rect 4351 2931 4387 2948
rect 4220 2891 4286 2907
rect 4220 2857 4236 2891
rect 4270 2857 4286 2891
rect 4328 2915 4394 2931
rect 4328 2881 4344 2915
rect 4378 2881 4394 2915
rect 4443 2907 4479 2948
rect 4328 2865 4394 2881
rect 4436 2891 4502 2907
rect 4220 2841 4286 2857
rect 4133 2819 4163 2834
rect 4251 2819 4281 2841
rect 4337 2819 4367 2865
rect 4436 2857 4452 2891
rect 4486 2857 4502 2891
rect 4436 2841 4502 2857
rect 4466 2819 4496 2841
rect 4544 2834 4580 2948
rect 4634 2931 4670 2948
rect 4753 2931 4789 2948
rect 4920 2946 4956 2963
rect 4622 2915 4688 2931
rect 4622 2881 4638 2915
rect 4672 2881 4688 2915
rect 4622 2865 4688 2881
rect 4736 2915 4802 2931
rect 4736 2881 4752 2915
rect 4786 2881 4802 2915
rect 4736 2868 4802 2881
rect 4920 2930 5054 2946
rect 4920 2896 4936 2930
rect 4970 2896 5004 2930
rect 5038 2896 5054 2930
rect 5171 2926 5207 2969
rect 5718 2967 5748 2982
rect 5821 2967 5851 2982
rect 5715 2940 5751 2967
rect 4920 2880 5054 2896
rect 5102 2910 5207 2926
rect 4544 2819 4574 2834
rect 4630 2819 4660 2865
rect 4736 2838 4872 2868
rect 4842 2819 4872 2838
rect 4987 2819 5017 2880
rect 5102 2876 5118 2910
rect 5152 2876 5207 2910
rect 5102 2860 5207 2876
rect 5703 2924 5769 2940
rect 5818 2924 5854 2967
rect 5919 2957 5955 2988
rect 6327 3161 6357 3187
rect 6428 3161 6458 3187
rect 6520 3161 6550 3187
rect 6618 3176 6654 3229
rect 6994 3191 7030 3229
rect 7248 3206 7278 3232
rect 6621 3161 6651 3176
rect 6711 3161 6741 3187
rect 6830 3161 6860 3187
rect 6997 3176 7027 3191
rect 7780 3202 7810 3228
rect 7981 3225 9092 3255
rect 7981 3214 8017 3225
rect 6997 2961 7027 2976
rect 7248 2967 7278 2982
rect 7883 3178 7913 3204
rect 7984 3199 8014 3214
rect 8085 3157 8115 3183
rect 8175 3157 8205 3183
rect 8269 3172 8305 3225
rect 8272 3157 8302 3172
rect 7984 2984 8014 2999
rect 5703 2890 5719 2924
rect 5753 2890 5769 2924
rect 5703 2874 5769 2890
rect 5811 2908 5877 2924
rect 5811 2874 5827 2908
rect 5861 2874 5877 2908
rect 5177 2838 5207 2860
rect 3644 2664 3674 2690
rect 3767 2665 3797 2691
rect 3845 2665 3875 2691
rect 3923 2665 3953 2691
rect 4031 2665 4061 2691
rect 4133 2665 4163 2691
rect 4251 2665 4281 2691
rect 4337 2665 4367 2691
rect 4466 2665 4496 2691
rect 4544 2665 4574 2691
rect 4630 2665 4660 2691
rect 4842 2665 4872 2691
rect 4987 2665 5017 2691
rect 5718 2836 5748 2874
rect 5811 2858 5877 2874
rect 5177 2664 5207 2690
rect 5841 2817 5871 2858
rect 5919 2817 5949 2957
rect 6023 2946 6053 2961
rect 6113 2946 6143 2961
rect 6210 2946 6240 2961
rect 6327 2946 6357 2961
rect 6428 2946 6458 2961
rect 6520 2946 6550 2961
rect 6621 2946 6651 2961
rect 6711 2946 6741 2961
rect 6830 2946 6860 2961
rect 6020 2929 6056 2946
rect 6110 2929 6146 2946
rect 5991 2913 6057 2929
rect 5991 2879 6007 2913
rect 6041 2879 6057 2913
rect 5991 2863 6057 2879
rect 6099 2913 6165 2929
rect 6099 2879 6115 2913
rect 6149 2879 6165 2913
rect 6099 2863 6165 2879
rect 5997 2817 6027 2863
rect 6105 2817 6135 2863
rect 6207 2832 6243 2946
rect 6324 2905 6360 2946
rect 6425 2929 6461 2946
rect 6294 2889 6360 2905
rect 6294 2855 6310 2889
rect 6344 2855 6360 2889
rect 6402 2913 6468 2929
rect 6402 2879 6418 2913
rect 6452 2879 6468 2913
rect 6517 2905 6553 2946
rect 6402 2863 6468 2879
rect 6510 2889 6576 2905
rect 6294 2839 6360 2855
rect 6207 2817 6237 2832
rect 6325 2817 6355 2839
rect 6411 2817 6441 2863
rect 6510 2855 6526 2889
rect 6560 2855 6576 2889
rect 6510 2839 6576 2855
rect 6540 2817 6570 2839
rect 6618 2832 6654 2946
rect 6708 2929 6744 2946
rect 6827 2929 6863 2946
rect 6994 2944 7030 2961
rect 6696 2913 6762 2929
rect 6696 2879 6712 2913
rect 6746 2879 6762 2913
rect 6696 2863 6762 2879
rect 6810 2913 6876 2929
rect 6810 2879 6826 2913
rect 6860 2879 6876 2913
rect 6810 2866 6876 2879
rect 6994 2928 7128 2944
rect 6994 2894 7010 2928
rect 7044 2894 7078 2928
rect 7112 2894 7128 2928
rect 7245 2924 7281 2967
rect 7780 2963 7810 2978
rect 7883 2963 7913 2978
rect 7777 2936 7813 2963
rect 6994 2878 7128 2894
rect 7176 2908 7281 2924
rect 6618 2817 6648 2832
rect 6704 2817 6734 2863
rect 6810 2836 6946 2866
rect 6916 2817 6946 2836
rect 7061 2817 7091 2878
rect 7176 2874 7192 2908
rect 7226 2874 7281 2908
rect 7176 2858 7281 2874
rect 7765 2920 7831 2936
rect 7880 2920 7916 2963
rect 7981 2953 8017 2984
rect 8389 3157 8419 3183
rect 8490 3157 8520 3183
rect 8582 3157 8612 3183
rect 8680 3172 8716 3225
rect 9056 3187 9092 3225
rect 9310 3202 9340 3228
rect 8683 3157 8713 3172
rect 8773 3157 8803 3183
rect 8892 3157 8922 3183
rect 9059 3172 9089 3187
rect 9840 3198 9870 3224
rect 10041 3221 11152 3251
rect 10041 3210 10077 3221
rect 9059 2957 9089 2972
rect 9310 2963 9340 2978
rect 9943 3174 9973 3200
rect 10044 3195 10074 3210
rect 10145 3153 10175 3179
rect 10235 3153 10265 3179
rect 10329 3168 10365 3221
rect 10332 3153 10362 3168
rect 10044 2980 10074 2995
rect 7765 2886 7781 2920
rect 7815 2886 7831 2920
rect 7765 2870 7831 2886
rect 7873 2904 7939 2920
rect 7873 2870 7889 2904
rect 7923 2870 7939 2904
rect 7251 2836 7281 2858
rect 5718 2662 5748 2688
rect 5841 2663 5871 2689
rect 5919 2663 5949 2689
rect 5997 2663 6027 2689
rect 6105 2663 6135 2689
rect 6207 2663 6237 2689
rect 6325 2663 6355 2689
rect 6411 2663 6441 2689
rect 6540 2663 6570 2689
rect 6618 2663 6648 2689
rect 6704 2663 6734 2689
rect 6916 2663 6946 2689
rect 7061 2663 7091 2689
rect 7780 2832 7810 2870
rect 7873 2854 7939 2870
rect 7251 2662 7281 2688
rect 7903 2813 7933 2854
rect 7981 2813 8011 2953
rect 8085 2942 8115 2957
rect 8175 2942 8205 2957
rect 8272 2942 8302 2957
rect 8389 2942 8419 2957
rect 8490 2942 8520 2957
rect 8582 2942 8612 2957
rect 8683 2942 8713 2957
rect 8773 2942 8803 2957
rect 8892 2942 8922 2957
rect 8082 2925 8118 2942
rect 8172 2925 8208 2942
rect 8053 2909 8119 2925
rect 8053 2875 8069 2909
rect 8103 2875 8119 2909
rect 8053 2859 8119 2875
rect 8161 2909 8227 2925
rect 8161 2875 8177 2909
rect 8211 2875 8227 2909
rect 8161 2859 8227 2875
rect 8059 2813 8089 2859
rect 8167 2813 8197 2859
rect 8269 2828 8305 2942
rect 8386 2901 8422 2942
rect 8487 2925 8523 2942
rect 8356 2885 8422 2901
rect 8356 2851 8372 2885
rect 8406 2851 8422 2885
rect 8464 2909 8530 2925
rect 8464 2875 8480 2909
rect 8514 2875 8530 2909
rect 8579 2901 8615 2942
rect 8464 2859 8530 2875
rect 8572 2885 8638 2901
rect 8356 2835 8422 2851
rect 8269 2813 8299 2828
rect 8387 2813 8417 2835
rect 8473 2813 8503 2859
rect 8572 2851 8588 2885
rect 8622 2851 8638 2885
rect 8572 2835 8638 2851
rect 8602 2813 8632 2835
rect 8680 2828 8716 2942
rect 8770 2925 8806 2942
rect 8889 2925 8925 2942
rect 9056 2940 9092 2957
rect 8758 2909 8824 2925
rect 8758 2875 8774 2909
rect 8808 2875 8824 2909
rect 8758 2859 8824 2875
rect 8872 2909 8938 2925
rect 8872 2875 8888 2909
rect 8922 2875 8938 2909
rect 8872 2862 8938 2875
rect 9056 2924 9190 2940
rect 9056 2890 9072 2924
rect 9106 2890 9140 2924
rect 9174 2890 9190 2924
rect 9307 2920 9343 2963
rect 9840 2959 9870 2974
rect 9943 2959 9973 2974
rect 9837 2932 9873 2959
rect 9056 2874 9190 2890
rect 9238 2904 9343 2920
rect 8680 2813 8710 2828
rect 8766 2813 8796 2859
rect 8872 2832 9008 2862
rect 8978 2813 9008 2832
rect 9123 2813 9153 2874
rect 9238 2870 9254 2904
rect 9288 2870 9343 2904
rect 9238 2854 9343 2870
rect 9825 2916 9891 2932
rect 9940 2916 9976 2959
rect 10041 2949 10077 2980
rect 10449 3153 10479 3179
rect 10550 3153 10580 3179
rect 10642 3153 10672 3179
rect 10740 3168 10776 3221
rect 11116 3183 11152 3221
rect 11370 3198 11400 3224
rect 10743 3153 10773 3168
rect 10833 3153 10863 3179
rect 10952 3153 10982 3179
rect 11119 3168 11149 3183
rect 11902 3194 11932 3220
rect 12103 3217 13214 3247
rect 12103 3206 12139 3217
rect 11119 2953 11149 2968
rect 11370 2959 11400 2974
rect 12005 3170 12035 3196
rect 12106 3191 12136 3206
rect 12207 3149 12237 3175
rect 12297 3149 12327 3175
rect 12391 3164 12427 3217
rect 12394 3149 12424 3164
rect 12106 2976 12136 2991
rect 9825 2882 9841 2916
rect 9875 2882 9891 2916
rect 9825 2866 9891 2882
rect 9933 2900 9999 2916
rect 9933 2866 9949 2900
rect 9983 2866 9999 2900
rect 9313 2832 9343 2854
rect 7780 2658 7810 2684
rect 7903 2659 7933 2685
rect 7981 2659 8011 2685
rect 8059 2659 8089 2685
rect 8167 2659 8197 2685
rect 8269 2659 8299 2685
rect 8387 2659 8417 2685
rect 8473 2659 8503 2685
rect 8602 2659 8632 2685
rect 8680 2659 8710 2685
rect 8766 2659 8796 2685
rect 8978 2659 9008 2685
rect 9123 2659 9153 2685
rect 9840 2828 9870 2866
rect 9933 2850 9999 2866
rect 9313 2658 9343 2684
rect 9963 2809 9993 2850
rect 10041 2809 10071 2949
rect 10145 2938 10175 2953
rect 10235 2938 10265 2953
rect 10332 2938 10362 2953
rect 10449 2938 10479 2953
rect 10550 2938 10580 2953
rect 10642 2938 10672 2953
rect 10743 2938 10773 2953
rect 10833 2938 10863 2953
rect 10952 2938 10982 2953
rect 10142 2921 10178 2938
rect 10232 2921 10268 2938
rect 10113 2905 10179 2921
rect 10113 2871 10129 2905
rect 10163 2871 10179 2905
rect 10113 2855 10179 2871
rect 10221 2905 10287 2921
rect 10221 2871 10237 2905
rect 10271 2871 10287 2905
rect 10221 2855 10287 2871
rect 10119 2809 10149 2855
rect 10227 2809 10257 2855
rect 10329 2824 10365 2938
rect 10446 2897 10482 2938
rect 10547 2921 10583 2938
rect 10416 2881 10482 2897
rect 10416 2847 10432 2881
rect 10466 2847 10482 2881
rect 10524 2905 10590 2921
rect 10524 2871 10540 2905
rect 10574 2871 10590 2905
rect 10639 2897 10675 2938
rect 10524 2855 10590 2871
rect 10632 2881 10698 2897
rect 10416 2831 10482 2847
rect 10329 2809 10359 2824
rect 10447 2809 10477 2831
rect 10533 2809 10563 2855
rect 10632 2847 10648 2881
rect 10682 2847 10698 2881
rect 10632 2831 10698 2847
rect 10662 2809 10692 2831
rect 10740 2824 10776 2938
rect 10830 2921 10866 2938
rect 10949 2921 10985 2938
rect 11116 2936 11152 2953
rect 10818 2905 10884 2921
rect 10818 2871 10834 2905
rect 10868 2871 10884 2905
rect 10818 2855 10884 2871
rect 10932 2905 10998 2921
rect 10932 2871 10948 2905
rect 10982 2871 10998 2905
rect 10932 2858 10998 2871
rect 11116 2920 11250 2936
rect 11116 2886 11132 2920
rect 11166 2886 11200 2920
rect 11234 2886 11250 2920
rect 11367 2916 11403 2959
rect 11902 2955 11932 2970
rect 12005 2955 12035 2970
rect 11899 2928 11935 2955
rect 11116 2870 11250 2886
rect 11298 2900 11403 2916
rect 10740 2809 10770 2824
rect 10826 2809 10856 2855
rect 10932 2828 11068 2858
rect 11038 2809 11068 2828
rect 11183 2809 11213 2870
rect 11298 2866 11314 2900
rect 11348 2866 11403 2900
rect 11298 2850 11403 2866
rect 11887 2912 11953 2928
rect 12002 2912 12038 2955
rect 12103 2945 12139 2976
rect 12511 3149 12541 3175
rect 12612 3149 12642 3175
rect 12704 3149 12734 3175
rect 12802 3164 12838 3217
rect 13178 3179 13214 3217
rect 13432 3194 13462 3220
rect 12805 3149 12835 3164
rect 12895 3149 12925 3175
rect 13014 3149 13044 3175
rect 13181 3164 13211 3179
rect 13976 3192 14006 3218
rect 14177 3215 15288 3245
rect 14177 3204 14213 3215
rect 13181 2949 13211 2964
rect 13432 2955 13462 2970
rect 14079 3168 14109 3194
rect 14180 3189 14210 3204
rect 14281 3147 14311 3173
rect 14371 3147 14401 3173
rect 14465 3162 14501 3215
rect 14468 3147 14498 3162
rect 14180 2974 14210 2989
rect 11887 2878 11903 2912
rect 11937 2878 11953 2912
rect 11887 2862 11953 2878
rect 11995 2896 12061 2912
rect 11995 2862 12011 2896
rect 12045 2862 12061 2896
rect 11373 2828 11403 2850
rect 9840 2654 9870 2680
rect 9963 2655 9993 2681
rect 10041 2655 10071 2681
rect 10119 2655 10149 2681
rect 10227 2655 10257 2681
rect 10329 2655 10359 2681
rect 10447 2655 10477 2681
rect 10533 2655 10563 2681
rect 10662 2655 10692 2681
rect 10740 2655 10770 2681
rect 10826 2655 10856 2681
rect 11038 2655 11068 2681
rect 11183 2655 11213 2681
rect 11902 2824 11932 2862
rect 11995 2846 12061 2862
rect 11373 2654 11403 2680
rect 12025 2805 12055 2846
rect 12103 2805 12133 2945
rect 12207 2934 12237 2949
rect 12297 2934 12327 2949
rect 12394 2934 12424 2949
rect 12511 2934 12541 2949
rect 12612 2934 12642 2949
rect 12704 2934 12734 2949
rect 12805 2934 12835 2949
rect 12895 2934 12925 2949
rect 13014 2934 13044 2949
rect 12204 2917 12240 2934
rect 12294 2917 12330 2934
rect 12175 2901 12241 2917
rect 12175 2867 12191 2901
rect 12225 2867 12241 2901
rect 12175 2851 12241 2867
rect 12283 2901 12349 2917
rect 12283 2867 12299 2901
rect 12333 2867 12349 2901
rect 12283 2851 12349 2867
rect 12181 2805 12211 2851
rect 12289 2805 12319 2851
rect 12391 2820 12427 2934
rect 12508 2893 12544 2934
rect 12609 2917 12645 2934
rect 12478 2877 12544 2893
rect 12478 2843 12494 2877
rect 12528 2843 12544 2877
rect 12586 2901 12652 2917
rect 12586 2867 12602 2901
rect 12636 2867 12652 2901
rect 12701 2893 12737 2934
rect 12586 2851 12652 2867
rect 12694 2877 12760 2893
rect 12478 2827 12544 2843
rect 12391 2805 12421 2820
rect 12509 2805 12539 2827
rect 12595 2805 12625 2851
rect 12694 2843 12710 2877
rect 12744 2843 12760 2877
rect 12694 2827 12760 2843
rect 12724 2805 12754 2827
rect 12802 2820 12838 2934
rect 12892 2917 12928 2934
rect 13011 2917 13047 2934
rect 13178 2932 13214 2949
rect 12880 2901 12946 2917
rect 12880 2867 12896 2901
rect 12930 2867 12946 2901
rect 12880 2851 12946 2867
rect 12994 2901 13060 2917
rect 12994 2867 13010 2901
rect 13044 2867 13060 2901
rect 12994 2854 13060 2867
rect 13178 2916 13312 2932
rect 13178 2882 13194 2916
rect 13228 2882 13262 2916
rect 13296 2882 13312 2916
rect 13429 2912 13465 2955
rect 13976 2953 14006 2968
rect 14079 2953 14109 2968
rect 13973 2926 14009 2953
rect 13178 2866 13312 2882
rect 13360 2896 13465 2912
rect 12802 2805 12832 2820
rect 12888 2805 12918 2851
rect 12994 2824 13130 2854
rect 13100 2805 13130 2824
rect 13245 2805 13275 2866
rect 13360 2862 13376 2896
rect 13410 2862 13465 2896
rect 13360 2846 13465 2862
rect 13961 2910 14027 2926
rect 14076 2910 14112 2953
rect 14177 2943 14213 2974
rect 14585 3147 14615 3173
rect 14686 3147 14716 3173
rect 14778 3147 14808 3173
rect 14876 3162 14912 3215
rect 15252 3177 15288 3215
rect 15506 3192 15536 3218
rect 14879 3147 14909 3162
rect 14969 3147 14999 3173
rect 15088 3147 15118 3173
rect 15255 3162 15285 3177
rect 16038 3188 16068 3214
rect 16239 3211 17350 3241
rect 16239 3200 16275 3211
rect 15255 2947 15285 2962
rect 15506 2953 15536 2968
rect 16141 3164 16171 3190
rect 16242 3185 16272 3200
rect 16343 3143 16373 3169
rect 16433 3143 16463 3169
rect 16527 3158 16563 3211
rect 16530 3143 16560 3158
rect 16242 2970 16272 2985
rect 13961 2876 13977 2910
rect 14011 2876 14027 2910
rect 13961 2860 14027 2876
rect 14069 2894 14135 2910
rect 14069 2860 14085 2894
rect 14119 2860 14135 2894
rect 13435 2824 13465 2846
rect 11902 2650 11932 2676
rect 12025 2651 12055 2677
rect 12103 2651 12133 2677
rect 12181 2651 12211 2677
rect 12289 2651 12319 2677
rect 12391 2651 12421 2677
rect 12509 2651 12539 2677
rect 12595 2651 12625 2677
rect 12724 2651 12754 2677
rect 12802 2651 12832 2677
rect 12888 2651 12918 2677
rect 13100 2651 13130 2677
rect 13245 2651 13275 2677
rect 13976 2822 14006 2860
rect 14069 2844 14135 2860
rect 13435 2650 13465 2676
rect 14099 2803 14129 2844
rect 14177 2803 14207 2943
rect 14281 2932 14311 2947
rect 14371 2932 14401 2947
rect 14468 2932 14498 2947
rect 14585 2932 14615 2947
rect 14686 2932 14716 2947
rect 14778 2932 14808 2947
rect 14879 2932 14909 2947
rect 14969 2932 14999 2947
rect 15088 2932 15118 2947
rect 14278 2915 14314 2932
rect 14368 2915 14404 2932
rect 14249 2899 14315 2915
rect 14249 2865 14265 2899
rect 14299 2865 14315 2899
rect 14249 2849 14315 2865
rect 14357 2899 14423 2915
rect 14357 2865 14373 2899
rect 14407 2865 14423 2899
rect 14357 2849 14423 2865
rect 14255 2803 14285 2849
rect 14363 2803 14393 2849
rect 14465 2818 14501 2932
rect 14582 2891 14618 2932
rect 14683 2915 14719 2932
rect 14552 2875 14618 2891
rect 14552 2841 14568 2875
rect 14602 2841 14618 2875
rect 14660 2899 14726 2915
rect 14660 2865 14676 2899
rect 14710 2865 14726 2899
rect 14775 2891 14811 2932
rect 14660 2849 14726 2865
rect 14768 2875 14834 2891
rect 14552 2825 14618 2841
rect 14465 2803 14495 2818
rect 14583 2803 14613 2825
rect 14669 2803 14699 2849
rect 14768 2841 14784 2875
rect 14818 2841 14834 2875
rect 14768 2825 14834 2841
rect 14798 2803 14828 2825
rect 14876 2818 14912 2932
rect 14966 2915 15002 2932
rect 15085 2915 15121 2932
rect 15252 2930 15288 2947
rect 14954 2899 15020 2915
rect 14954 2865 14970 2899
rect 15004 2865 15020 2899
rect 14954 2849 15020 2865
rect 15068 2899 15134 2915
rect 15068 2865 15084 2899
rect 15118 2865 15134 2899
rect 15068 2852 15134 2865
rect 15252 2914 15386 2930
rect 15252 2880 15268 2914
rect 15302 2880 15336 2914
rect 15370 2880 15386 2914
rect 15503 2910 15539 2953
rect 16038 2949 16068 2964
rect 16141 2949 16171 2964
rect 16035 2922 16071 2949
rect 15252 2864 15386 2880
rect 15434 2894 15539 2910
rect 14876 2803 14906 2818
rect 14962 2803 14992 2849
rect 15068 2822 15204 2852
rect 15174 2803 15204 2822
rect 15319 2803 15349 2864
rect 15434 2860 15450 2894
rect 15484 2860 15539 2894
rect 15434 2844 15539 2860
rect 16023 2906 16089 2922
rect 16138 2906 16174 2949
rect 16239 2939 16275 2970
rect 16647 3143 16677 3169
rect 16748 3143 16778 3169
rect 16840 3143 16870 3169
rect 16938 3158 16974 3211
rect 17314 3173 17350 3211
rect 17568 3188 17598 3214
rect 16941 3143 16971 3158
rect 17031 3143 17061 3169
rect 17150 3143 17180 3169
rect 17317 3158 17347 3173
rect 22664 3083 22694 3109
rect 17317 2943 17347 2958
rect 17568 2949 17598 2964
rect 16023 2872 16039 2906
rect 16073 2872 16089 2906
rect 16023 2856 16089 2872
rect 16131 2890 16197 2906
rect 16131 2856 16147 2890
rect 16181 2856 16197 2890
rect 15509 2822 15539 2844
rect 13976 2648 14006 2674
rect 14099 2649 14129 2675
rect 14177 2649 14207 2675
rect 14255 2649 14285 2675
rect 14363 2649 14393 2675
rect 14465 2649 14495 2675
rect 14583 2649 14613 2675
rect 14669 2649 14699 2675
rect 14798 2649 14828 2675
rect 14876 2649 14906 2675
rect 14962 2649 14992 2675
rect 15174 2649 15204 2675
rect 15319 2649 15349 2675
rect 16038 2818 16068 2856
rect 16131 2840 16197 2856
rect 15509 2648 15539 2674
rect 16161 2799 16191 2840
rect 16239 2799 16269 2939
rect 16343 2928 16373 2943
rect 16433 2928 16463 2943
rect 16530 2928 16560 2943
rect 16647 2928 16677 2943
rect 16748 2928 16778 2943
rect 16840 2928 16870 2943
rect 16941 2928 16971 2943
rect 17031 2928 17061 2943
rect 17150 2928 17180 2943
rect 16340 2911 16376 2928
rect 16430 2911 16466 2928
rect 16311 2895 16377 2911
rect 16311 2861 16327 2895
rect 16361 2861 16377 2895
rect 16311 2845 16377 2861
rect 16419 2895 16485 2911
rect 16419 2861 16435 2895
rect 16469 2861 16485 2895
rect 16419 2845 16485 2861
rect 16317 2799 16347 2845
rect 16425 2799 16455 2845
rect 16527 2814 16563 2928
rect 16644 2887 16680 2928
rect 16745 2911 16781 2928
rect 16614 2871 16680 2887
rect 16614 2837 16630 2871
rect 16664 2837 16680 2871
rect 16722 2895 16788 2911
rect 16722 2861 16738 2895
rect 16772 2861 16788 2895
rect 16837 2887 16873 2928
rect 16722 2845 16788 2861
rect 16830 2871 16896 2887
rect 16614 2821 16680 2837
rect 16527 2799 16557 2814
rect 16645 2799 16675 2821
rect 16731 2799 16761 2845
rect 16830 2837 16846 2871
rect 16880 2837 16896 2871
rect 16830 2821 16896 2837
rect 16860 2799 16890 2821
rect 16938 2814 16974 2928
rect 17028 2911 17064 2928
rect 17147 2911 17183 2928
rect 17314 2926 17350 2943
rect 17016 2895 17082 2911
rect 17016 2861 17032 2895
rect 17066 2861 17082 2895
rect 17016 2845 17082 2861
rect 17130 2895 17196 2911
rect 17130 2861 17146 2895
rect 17180 2861 17196 2895
rect 17130 2848 17196 2861
rect 17314 2910 17448 2926
rect 17314 2876 17330 2910
rect 17364 2876 17398 2910
rect 17432 2876 17448 2910
rect 17565 2906 17601 2949
rect 17314 2860 17448 2876
rect 17496 2890 17601 2906
rect 16938 2799 16968 2814
rect 17024 2799 17054 2845
rect 17130 2818 17266 2848
rect 17236 2799 17266 2818
rect 17381 2799 17411 2860
rect 17496 2856 17512 2890
rect 17546 2856 17601 2890
rect 23249 3081 23279 3107
rect 23333 3081 23363 3107
rect 17496 2840 17601 2856
rect 22664 2851 22694 2883
rect 23865 3069 23895 3095
rect 23949 3069 23979 3095
rect 24033 3069 24063 3095
rect 24117 3069 24147 3095
rect 17571 2818 17601 2840
rect 22608 2835 22694 2851
rect 23249 2849 23279 2881
rect 23333 2849 23363 2881
rect 24713 3055 24743 3081
rect 24797 3055 24827 3081
rect 24881 3055 24911 3081
rect 24965 3055 24995 3081
rect 25049 3055 25079 3081
rect 25133 3055 25163 3081
rect 16038 2644 16068 2670
rect 16161 2645 16191 2671
rect 16239 2645 16269 2671
rect 16317 2645 16347 2671
rect 16425 2645 16455 2671
rect 16527 2645 16557 2671
rect 16645 2645 16675 2671
rect 16731 2645 16761 2671
rect 16860 2645 16890 2671
rect 16938 2645 16968 2671
rect 17024 2645 17054 2671
rect 17236 2645 17266 2671
rect 17381 2645 17411 2671
rect 22608 2801 22624 2835
rect 22658 2801 22694 2835
rect 22608 2785 22694 2801
rect 22664 2763 22694 2785
rect 23189 2833 23363 2849
rect 23865 2837 23895 2869
rect 23949 2837 23979 2869
rect 24033 2837 24063 2869
rect 24117 2837 24147 2869
rect 23189 2799 23205 2833
rect 23239 2799 23363 2833
rect 23189 2783 23363 2799
rect 17571 2644 17601 2670
rect 23249 2761 23279 2783
rect 23333 2761 23363 2783
rect 23797 2821 24147 2837
rect 24713 2823 24743 2855
rect 24797 2823 24827 2855
rect 24881 2823 24911 2855
rect 24965 2823 24995 2855
rect 25049 2823 25079 2855
rect 25133 2823 25163 2855
rect 23797 2787 23813 2821
rect 23847 2787 23905 2821
rect 23939 2787 23989 2821
rect 24023 2787 24073 2821
rect 24107 2787 24147 2821
rect 23797 2771 24147 2787
rect 22664 2607 22694 2633
rect 23865 2749 23895 2771
rect 23949 2749 23979 2771
rect 24033 2749 24063 2771
rect 24117 2749 24147 2771
rect 24621 2807 25163 2823
rect 24621 2773 24637 2807
rect 24671 2773 24905 2807
rect 24939 2773 24989 2807
rect 25023 2773 25073 2807
rect 25107 2773 25163 2807
rect 24621 2757 25163 2773
rect 23249 2605 23279 2631
rect 23333 2605 23363 2631
rect 24713 2735 24743 2757
rect 24797 2735 24827 2757
rect 24881 2735 24911 2757
rect 24965 2735 24995 2757
rect 25049 2735 25079 2757
rect 25133 2735 25163 2757
rect 23865 2593 23895 2619
rect 23949 2593 23979 2619
rect 24033 2593 24063 2619
rect 24117 2593 24147 2619
rect 24713 2579 24743 2605
rect 24797 2579 24827 2605
rect 24881 2579 24911 2605
rect 24965 2579 24995 2605
rect 25049 2579 25079 2605
rect 25133 2579 25163 2605
<< polycont >>
rect 8315 4142 8349 4176
rect 1583 2896 1617 2930
rect 1691 2880 1725 2914
rect 1871 2885 1905 2919
rect 1979 2885 2013 2919
rect 2174 2861 2208 2895
rect 2282 2885 2316 2919
rect 2390 2861 2424 2895
rect 2576 2885 2610 2919
rect 2690 2885 2724 2919
rect 2874 2900 2908 2934
rect 2942 2900 2976 2934
rect 3056 2880 3090 2914
rect 3645 2892 3679 2926
rect 3753 2876 3787 2910
rect 3933 2881 3967 2915
rect 4041 2881 4075 2915
rect 4236 2857 4270 2891
rect 4344 2881 4378 2915
rect 4452 2857 4486 2891
rect 4638 2881 4672 2915
rect 4752 2881 4786 2915
rect 4936 2896 4970 2930
rect 5004 2896 5038 2930
rect 5118 2876 5152 2910
rect 5719 2890 5753 2924
rect 5827 2874 5861 2908
rect 6007 2879 6041 2913
rect 6115 2879 6149 2913
rect 6310 2855 6344 2889
rect 6418 2879 6452 2913
rect 6526 2855 6560 2889
rect 6712 2879 6746 2913
rect 6826 2879 6860 2913
rect 7010 2894 7044 2928
rect 7078 2894 7112 2928
rect 7192 2874 7226 2908
rect 7781 2886 7815 2920
rect 7889 2870 7923 2904
rect 8069 2875 8103 2909
rect 8177 2875 8211 2909
rect 8372 2851 8406 2885
rect 8480 2875 8514 2909
rect 8588 2851 8622 2885
rect 8774 2875 8808 2909
rect 8888 2875 8922 2909
rect 9072 2890 9106 2924
rect 9140 2890 9174 2924
rect 9254 2870 9288 2904
rect 9841 2882 9875 2916
rect 9949 2866 9983 2900
rect 10129 2871 10163 2905
rect 10237 2871 10271 2905
rect 10432 2847 10466 2881
rect 10540 2871 10574 2905
rect 10648 2847 10682 2881
rect 10834 2871 10868 2905
rect 10948 2871 10982 2905
rect 11132 2886 11166 2920
rect 11200 2886 11234 2920
rect 11314 2866 11348 2900
rect 11903 2878 11937 2912
rect 12011 2862 12045 2896
rect 12191 2867 12225 2901
rect 12299 2867 12333 2901
rect 12494 2843 12528 2877
rect 12602 2867 12636 2901
rect 12710 2843 12744 2877
rect 12896 2867 12930 2901
rect 13010 2867 13044 2901
rect 13194 2882 13228 2916
rect 13262 2882 13296 2916
rect 13376 2862 13410 2896
rect 13977 2876 14011 2910
rect 14085 2860 14119 2894
rect 14265 2865 14299 2899
rect 14373 2865 14407 2899
rect 14568 2841 14602 2875
rect 14676 2865 14710 2899
rect 14784 2841 14818 2875
rect 14970 2865 15004 2899
rect 15084 2865 15118 2899
rect 15268 2880 15302 2914
rect 15336 2880 15370 2914
rect 15450 2860 15484 2894
rect 16039 2872 16073 2906
rect 16147 2856 16181 2890
rect 16327 2861 16361 2895
rect 16435 2861 16469 2895
rect 16630 2837 16664 2871
rect 16738 2861 16772 2895
rect 16846 2837 16880 2871
rect 17032 2861 17066 2895
rect 17146 2861 17180 2895
rect 17330 2876 17364 2910
rect 17398 2876 17432 2910
rect 17512 2856 17546 2890
rect 22624 2801 22658 2835
rect 23205 2799 23239 2833
rect 23813 2787 23847 2821
rect 23905 2787 23939 2821
rect 23989 2787 24023 2821
rect 24073 2787 24107 2821
rect 24637 2773 24671 2807
rect 24905 2773 24939 2807
rect 24989 2773 25023 2807
rect 25073 2773 25107 2807
<< locali >>
rect 8098 4435 8129 4469
rect 8163 4435 8225 4469
rect 8259 4435 8321 4469
rect 8355 4435 8386 4469
rect 8122 4366 8172 4435
rect 8122 4332 8138 4366
rect 8122 4276 8172 4332
rect 8122 4242 8138 4276
rect 8122 4226 8172 4242
rect 8208 4366 8274 4382
rect 8208 4332 8224 4366
rect 8258 4332 8274 4366
rect 8208 4276 8274 4332
rect 8208 4242 8224 4276
rect 8258 4242 8274 4276
rect 8208 4226 8274 4242
rect 8310 4366 8360 4435
rect 8344 4332 8360 4366
rect 8310 4276 8360 4332
rect 8344 4242 8360 4276
rect 8310 4226 8360 4242
rect 8208 4138 8265 4226
rect 8208 4096 8220 4138
rect 8256 4096 8265 4138
rect 8299 4176 8365 4192
rect 8299 4142 8315 4176
rect 8349 4146 8365 4176
rect 8299 4112 8320 4142
rect 8354 4112 8365 4146
rect 8299 4096 8365 4112
rect 8119 4072 8169 4088
rect 8119 4038 8135 4072
rect 8119 3989 8169 4038
rect 8119 3955 8135 3989
rect 8119 3906 8169 3955
rect 8119 3872 8135 3906
rect 8119 3803 8169 3872
rect 8208 4072 8265 4096
rect 8208 4038 8225 4072
rect 8259 4038 8265 4072
rect 8208 3989 8265 4038
rect 8208 3955 8225 3989
rect 8259 3955 8265 3989
rect 8208 3906 8265 3955
rect 8208 3872 8225 3906
rect 8259 3872 8265 3906
rect 8208 3856 8265 3872
rect 8299 4046 8365 4062
rect 8299 4012 8315 4046
rect 8349 4012 8365 4046
rect 8299 3976 8365 4012
rect 8299 3942 8315 3976
rect 8349 3942 8365 3976
rect 8299 3906 8365 3942
rect 8299 3872 8315 3906
rect 8349 3872 8365 3906
rect 8299 3803 8365 3872
rect 8098 3769 8129 3803
rect 8163 3769 8225 3803
rect 8259 3769 8321 3803
rect 8355 3769 8386 3803
rect 1498 3269 1529 3303
rect 1563 3269 1625 3303
rect 1659 3269 1721 3303
rect 1755 3269 1817 3303
rect 1851 3269 1913 3303
rect 1947 3269 2009 3303
rect 2043 3269 2105 3303
rect 2139 3269 2201 3303
rect 2235 3269 2297 3303
rect 2331 3269 2393 3303
rect 2427 3269 2489 3303
rect 2523 3269 2585 3303
rect 2619 3269 2681 3303
rect 2715 3269 2777 3303
rect 2811 3269 2873 3303
rect 2907 3269 2969 3303
rect 3003 3269 3065 3303
rect 3099 3269 3161 3303
rect 3195 3269 3226 3303
rect 1515 3200 1569 3216
rect 1515 3166 1535 3200
rect 1515 3117 1569 3166
rect 1515 3083 1535 3117
rect 1515 3034 1569 3083
rect 1515 3000 1535 3034
rect 1609 3200 1675 3269
rect 1609 3166 1625 3200
rect 1659 3166 1675 3200
rect 2114 3196 2180 3269
rect 1609 3132 1675 3166
rect 1609 3098 1625 3132
rect 1659 3098 1675 3132
rect 1609 3064 1675 3098
rect 1609 3030 1625 3064
rect 1659 3030 1675 3064
rect 1914 3155 1980 3171
rect 1914 3121 1930 3155
rect 1964 3121 1980 3155
rect 1914 3087 1980 3121
rect 1914 3053 1930 3087
rect 1964 3053 1980 3087
rect 1914 3044 1980 3053
rect 1515 2984 1569 3000
rect 1709 3019 1980 3044
rect 1709 3010 1930 3019
rect 1709 2996 1743 3010
rect 1515 2846 1549 2984
rect 1605 2962 1743 2996
rect 1914 2985 1930 3010
rect 1964 2985 1980 3019
rect 2020 3155 2070 3171
rect 2054 3121 2070 3155
rect 2114 3162 2130 3196
rect 2164 3162 2180 3196
rect 2114 3146 2180 3162
rect 2020 3112 2070 3121
rect 2218 3128 2284 3171
rect 2218 3112 2234 3128
rect 2020 3094 2234 3112
rect 2268 3094 2284 3128
rect 2020 3078 2284 3094
rect 2319 3131 2385 3269
rect 2319 3097 2335 3131
rect 2369 3097 2385 3131
rect 2319 3081 2385 3097
rect 2512 3155 2597 3171
rect 2512 3121 2528 3155
rect 2562 3121 2597 3155
rect 2020 3063 2070 3078
rect 2054 3029 2070 3063
rect 2512 3044 2597 3121
rect 2020 3013 2070 3029
rect 1811 2970 1857 2976
rect 1605 2946 1639 2962
rect 1583 2930 1639 2946
rect 1617 2896 1639 2930
rect 1811 2936 1817 2970
rect 1851 2936 1857 2970
rect 1914 2969 1980 2985
rect 2104 3010 2528 3044
rect 2562 3010 2597 3044
rect 2631 3155 2688 3171
rect 2631 3121 2647 3155
rect 2681 3121 2688 3155
rect 2631 3071 2688 3121
rect 2722 3157 2863 3269
rect 3049 3200 3115 3269
rect 3560 3265 3591 3299
rect 3625 3265 3687 3299
rect 3721 3265 3783 3299
rect 3817 3265 3879 3299
rect 3913 3265 3975 3299
rect 4009 3265 4071 3299
rect 4105 3265 4167 3299
rect 4201 3265 4263 3299
rect 4297 3265 4359 3299
rect 4393 3265 4455 3299
rect 4489 3265 4551 3299
rect 4585 3265 4647 3299
rect 4681 3265 4743 3299
rect 4777 3265 4839 3299
rect 4873 3265 4935 3299
rect 4969 3265 5031 3299
rect 5065 3265 5127 3299
rect 5161 3265 5223 3299
rect 5257 3265 5288 3299
rect 2722 3123 2738 3157
rect 2772 3123 2813 3157
rect 2847 3123 2863 3157
rect 2722 3120 2863 3123
rect 2898 3170 2962 3186
rect 2898 3136 2912 3170
rect 2946 3136 2962 3170
rect 2898 3071 2962 3136
rect 2631 3037 2647 3071
rect 2681 3060 2962 3071
rect 2681 3037 2912 3060
rect 2896 3026 2912 3037
rect 2946 3026 2962 3060
rect 2896 3010 2962 3026
rect 3049 3166 3065 3200
rect 3099 3166 3115 3200
rect 3049 3117 3115 3166
rect 3049 3083 3065 3117
rect 3099 3083 3115 3117
rect 3049 3034 3115 3083
rect 2104 2979 2138 3010
rect 1811 2935 1857 2936
rect 2014 2945 2138 2979
rect 2563 3003 2597 3010
rect 2266 2970 2337 2976
rect 2014 2935 2048 2945
rect 1583 2880 1639 2896
rect 1515 2830 1571 2846
rect 1515 2796 1537 2830
rect 1515 2740 1571 2796
rect 1515 2706 1537 2740
rect 1605 2770 1639 2880
rect 1675 2914 1741 2928
rect 1675 2880 1691 2914
rect 1725 2880 1741 2914
rect 1675 2864 1741 2880
rect 1811 2919 1921 2935
rect 1811 2885 1871 2919
rect 1905 2885 1921 2919
rect 1811 2872 1921 2885
rect 1963 2919 2048 2935
rect 1963 2885 1979 2919
rect 2013 2885 2048 2919
rect 2266 2936 2297 2970
rect 2331 2936 2337 2970
rect 2266 2919 2337 2936
rect 1963 2872 2048 2885
rect 2158 2895 2224 2911
rect 1707 2838 1741 2864
rect 2158 2861 2174 2895
rect 2208 2861 2224 2895
rect 2266 2885 2282 2919
rect 2316 2885 2337 2919
rect 2483 2970 2529 2976
rect 2483 2936 2489 2970
rect 2523 2936 2529 2970
rect 2563 2969 2808 3003
rect 3049 3000 3065 3034
rect 3099 3000 3115 3034
rect 3049 2984 3115 3000
rect 3155 3200 3206 3216
rect 3189 3166 3206 3200
rect 3155 3117 3206 3166
rect 3189 3083 3206 3117
rect 3155 3034 3206 3083
rect 3189 3000 3206 3034
rect 2483 2935 2529 2936
rect 2483 2919 2626 2935
rect 2266 2872 2337 2885
rect 2374 2896 2440 2911
rect 2374 2895 2396 2896
rect 2158 2838 2224 2861
rect 2374 2861 2390 2895
rect 2430 2862 2440 2896
rect 2483 2885 2576 2919
rect 2610 2885 2626 2919
rect 2483 2875 2626 2885
rect 2660 2919 2740 2935
rect 2660 2885 2690 2919
rect 2724 2885 2740 2919
rect 2660 2884 2740 2885
rect 2424 2861 2440 2862
rect 2374 2841 2440 2861
rect 2660 2841 2694 2884
rect 2774 2850 2808 2969
rect 2858 2940 2992 2976
rect 2858 2934 2920 2940
rect 2960 2934 2992 2940
rect 2858 2900 2874 2934
rect 2908 2900 2920 2934
rect 2976 2900 2992 2934
rect 3155 2960 3206 3000
rect 3577 3196 3631 3212
rect 3577 3162 3597 3196
rect 3577 3113 3631 3162
rect 3577 3079 3597 3113
rect 3577 3030 3631 3079
rect 3577 2996 3597 3030
rect 3671 3196 3737 3265
rect 3671 3162 3687 3196
rect 3721 3162 3737 3196
rect 4176 3192 4242 3265
rect 3671 3128 3737 3162
rect 3671 3094 3687 3128
rect 3721 3094 3737 3128
rect 3671 3060 3737 3094
rect 3671 3026 3687 3060
rect 3721 3026 3737 3060
rect 3976 3151 4042 3167
rect 3976 3117 3992 3151
rect 4026 3117 4042 3151
rect 3976 3083 4042 3117
rect 3976 3049 3992 3083
rect 4026 3049 4042 3083
rect 3976 3040 4042 3049
rect 3577 2980 3631 2996
rect 3771 3015 4042 3040
rect 3771 3006 3992 3015
rect 3771 2992 3805 3006
rect 2858 2898 2920 2900
rect 2960 2898 2992 2900
rect 2858 2884 2992 2898
rect 3040 2914 3106 2930
rect 3040 2880 3056 2914
rect 3090 2880 3106 2914
rect 3040 2850 3106 2880
rect 2374 2838 2694 2841
rect 1707 2807 2694 2838
rect 2728 2816 3106 2850
rect 3155 2926 3174 2960
rect 3155 2846 3206 2926
rect 3140 2830 3206 2846
rect 1707 2804 2440 2807
rect 2728 2773 2762 2816
rect 3140 2796 3156 2830
rect 3190 2796 3206 2830
rect 1605 2747 1952 2770
rect 1605 2736 1902 2747
rect 1515 2690 1571 2706
rect 1886 2713 1902 2736
rect 1936 2713 1952 2747
rect 1623 2668 1641 2702
rect 1675 2668 1694 2702
rect 1886 2691 1952 2713
rect 1994 2754 2280 2770
rect 1994 2720 2018 2754
rect 2052 2736 2230 2754
rect 2052 2720 2076 2736
rect 1994 2704 2076 2720
rect 2214 2720 2230 2736
rect 2264 2720 2280 2754
rect 2214 2704 2280 2720
rect 2314 2746 2409 2762
rect 2314 2712 2344 2746
rect 2378 2712 2409 2746
rect 1623 2637 1694 2668
rect 2112 2668 2128 2702
rect 2162 2668 2178 2702
rect 2112 2637 2178 2668
rect 2314 2637 2409 2712
rect 2507 2757 2762 2773
rect 2507 2723 2523 2757
rect 2557 2739 2762 2757
rect 2796 2766 3016 2782
rect 2796 2748 2966 2766
rect 2557 2723 2573 2739
rect 2507 2707 2573 2723
rect 2796 2705 2830 2748
rect 2950 2732 2966 2748
rect 3000 2732 3016 2766
rect 2950 2716 3016 2732
rect 3054 2758 3104 2774
rect 3054 2724 3070 2758
rect 2609 2671 2625 2705
rect 2659 2671 2719 2705
rect 2753 2671 2830 2705
rect 2864 2698 2914 2714
rect 2898 2664 2914 2698
rect 2864 2637 2914 2664
rect 3054 2637 3104 2724
rect 3140 2740 3206 2796
rect 3140 2706 3156 2740
rect 3190 2706 3206 2740
rect 3140 2690 3206 2706
rect 3577 2842 3611 2980
rect 3667 2958 3805 2992
rect 3976 2981 3992 3006
rect 4026 2981 4042 3015
rect 4082 3151 4132 3167
rect 4116 3117 4132 3151
rect 4176 3158 4192 3192
rect 4226 3158 4242 3192
rect 4176 3142 4242 3158
rect 4082 3108 4132 3117
rect 4280 3124 4346 3167
rect 4280 3108 4296 3124
rect 4082 3090 4296 3108
rect 4330 3090 4346 3124
rect 4082 3074 4346 3090
rect 4381 3127 4447 3265
rect 4381 3093 4397 3127
rect 4431 3093 4447 3127
rect 4381 3077 4447 3093
rect 4574 3151 4659 3167
rect 4574 3117 4590 3151
rect 4624 3117 4659 3151
rect 4082 3059 4132 3074
rect 4116 3025 4132 3059
rect 4574 3040 4659 3117
rect 4082 3009 4132 3025
rect 3873 2966 3919 2972
rect 3667 2942 3701 2958
rect 3645 2926 3701 2942
rect 3679 2892 3701 2926
rect 3873 2932 3879 2966
rect 3913 2932 3919 2966
rect 3976 2965 4042 2981
rect 4166 3006 4590 3040
rect 4624 3006 4659 3040
rect 4693 3151 4750 3167
rect 4693 3117 4709 3151
rect 4743 3117 4750 3151
rect 4693 3067 4750 3117
rect 4784 3153 4925 3265
rect 5111 3196 5177 3265
rect 5634 3263 5665 3297
rect 5699 3263 5761 3297
rect 5795 3263 5857 3297
rect 5891 3263 5953 3297
rect 5987 3263 6049 3297
rect 6083 3263 6145 3297
rect 6179 3263 6241 3297
rect 6275 3263 6337 3297
rect 6371 3263 6433 3297
rect 6467 3263 6529 3297
rect 6563 3263 6625 3297
rect 6659 3263 6721 3297
rect 6755 3263 6817 3297
rect 6851 3263 6913 3297
rect 6947 3263 7009 3297
rect 7043 3263 7105 3297
rect 7139 3263 7201 3297
rect 7235 3263 7297 3297
rect 7331 3263 7362 3297
rect 4784 3119 4800 3153
rect 4834 3119 4875 3153
rect 4909 3119 4925 3153
rect 4784 3116 4925 3119
rect 4960 3166 5024 3182
rect 4960 3132 4974 3166
rect 5008 3132 5024 3166
rect 4960 3067 5024 3132
rect 4693 3033 4709 3067
rect 4743 3056 5024 3067
rect 4743 3033 4974 3056
rect 4958 3022 4974 3033
rect 5008 3022 5024 3056
rect 4958 3006 5024 3022
rect 5111 3162 5127 3196
rect 5161 3162 5177 3196
rect 5111 3113 5177 3162
rect 5111 3079 5127 3113
rect 5161 3079 5177 3113
rect 5111 3030 5177 3079
rect 4166 2975 4200 3006
rect 3873 2931 3919 2932
rect 4076 2941 4200 2975
rect 4625 2999 4659 3006
rect 4328 2966 4399 2972
rect 4076 2931 4110 2941
rect 3645 2876 3701 2892
rect 3577 2826 3633 2842
rect 3577 2792 3599 2826
rect 3577 2736 3633 2792
rect 3577 2702 3599 2736
rect 3667 2766 3701 2876
rect 3737 2910 3803 2924
rect 3737 2876 3753 2910
rect 3787 2876 3803 2910
rect 3737 2860 3803 2876
rect 3873 2915 3983 2931
rect 3873 2881 3933 2915
rect 3967 2881 3983 2915
rect 3873 2868 3983 2881
rect 4025 2915 4110 2931
rect 4025 2881 4041 2915
rect 4075 2881 4110 2915
rect 4328 2932 4359 2966
rect 4393 2932 4399 2966
rect 4328 2915 4399 2932
rect 4025 2868 4110 2881
rect 4220 2891 4286 2907
rect 3769 2834 3803 2860
rect 4220 2857 4236 2891
rect 4270 2857 4286 2891
rect 4328 2881 4344 2915
rect 4378 2881 4399 2915
rect 4545 2966 4591 2972
rect 4545 2932 4551 2966
rect 4585 2932 4591 2966
rect 4625 2965 4870 2999
rect 5111 2996 5127 3030
rect 5161 2996 5177 3030
rect 5111 2980 5177 2996
rect 5217 3196 5268 3212
rect 5251 3162 5268 3196
rect 5217 3113 5268 3162
rect 5251 3079 5268 3113
rect 5217 3030 5268 3079
rect 5251 2996 5268 3030
rect 4545 2931 4591 2932
rect 4545 2915 4688 2931
rect 4328 2868 4399 2881
rect 4436 2892 4502 2907
rect 4436 2891 4458 2892
rect 4220 2834 4286 2857
rect 4436 2857 4452 2891
rect 4492 2858 4502 2892
rect 4545 2881 4638 2915
rect 4672 2881 4688 2915
rect 4545 2871 4688 2881
rect 4722 2915 4802 2931
rect 4722 2881 4752 2915
rect 4786 2881 4802 2915
rect 4722 2880 4802 2881
rect 4486 2857 4502 2858
rect 4436 2837 4502 2857
rect 4722 2837 4756 2880
rect 4836 2846 4870 2965
rect 4920 2936 5054 2972
rect 4920 2930 4982 2936
rect 5022 2930 5054 2936
rect 4920 2896 4936 2930
rect 4970 2896 4982 2930
rect 5038 2896 5054 2930
rect 5217 2962 5268 2996
rect 5217 2928 5232 2962
rect 4920 2894 4982 2896
rect 5022 2894 5054 2896
rect 4920 2880 5054 2894
rect 5102 2910 5168 2926
rect 5102 2876 5118 2910
rect 5152 2876 5168 2910
rect 5102 2846 5168 2876
rect 4436 2834 4756 2837
rect 3769 2803 4756 2834
rect 4790 2812 5168 2846
rect 5217 2842 5268 2928
rect 5202 2826 5268 2842
rect 3769 2800 4502 2803
rect 4790 2769 4824 2812
rect 5202 2792 5218 2826
rect 5252 2792 5268 2826
rect 3667 2743 4014 2766
rect 3667 2732 3964 2743
rect 3577 2686 3633 2702
rect 3948 2709 3964 2732
rect 3998 2709 4014 2743
rect 3685 2664 3703 2698
rect 3737 2664 3756 2698
rect 3948 2687 4014 2709
rect 4056 2750 4342 2766
rect 4056 2716 4080 2750
rect 4114 2732 4292 2750
rect 4114 2716 4138 2732
rect 4056 2700 4138 2716
rect 4276 2716 4292 2732
rect 4326 2716 4342 2750
rect 4276 2700 4342 2716
rect 4376 2742 4471 2758
rect 4376 2708 4406 2742
rect 4440 2708 4471 2742
rect 1498 2603 1529 2637
rect 1563 2603 1625 2637
rect 1659 2603 1721 2637
rect 1755 2603 1817 2637
rect 1851 2603 1913 2637
rect 1947 2603 2009 2637
rect 2043 2603 2105 2637
rect 2139 2603 2201 2637
rect 2235 2603 2297 2637
rect 2331 2603 2393 2637
rect 2427 2603 2489 2637
rect 2523 2603 2585 2637
rect 2619 2603 2681 2637
rect 2715 2603 2777 2637
rect 2811 2603 2873 2637
rect 2907 2603 2969 2637
rect 3003 2603 3065 2637
rect 3099 2603 3161 2637
rect 3195 2603 3226 2637
rect 3685 2633 3756 2664
rect 4174 2664 4190 2698
rect 4224 2664 4240 2698
rect 4174 2633 4240 2664
rect 4376 2633 4471 2708
rect 4569 2753 4824 2769
rect 4569 2719 4585 2753
rect 4619 2735 4824 2753
rect 4858 2762 5078 2778
rect 4858 2744 5028 2762
rect 4619 2719 4635 2735
rect 4569 2703 4635 2719
rect 4858 2701 4892 2744
rect 5012 2728 5028 2744
rect 5062 2728 5078 2762
rect 5012 2712 5078 2728
rect 5116 2754 5166 2770
rect 5116 2720 5132 2754
rect 4671 2667 4687 2701
rect 4721 2667 4781 2701
rect 4815 2667 4892 2701
rect 4926 2694 4976 2710
rect 4960 2660 4976 2694
rect 4926 2633 4976 2660
rect 5116 2633 5166 2720
rect 5202 2736 5268 2792
rect 5202 2702 5218 2736
rect 5252 2702 5268 2736
rect 5202 2686 5268 2702
rect 5651 3194 5705 3210
rect 5651 3160 5671 3194
rect 5651 3111 5705 3160
rect 5651 3077 5671 3111
rect 5651 3028 5705 3077
rect 5651 2994 5671 3028
rect 5745 3194 5811 3263
rect 5745 3160 5761 3194
rect 5795 3160 5811 3194
rect 6250 3190 6316 3263
rect 5745 3126 5811 3160
rect 5745 3092 5761 3126
rect 5795 3092 5811 3126
rect 5745 3058 5811 3092
rect 5745 3024 5761 3058
rect 5795 3024 5811 3058
rect 6050 3149 6116 3165
rect 6050 3115 6066 3149
rect 6100 3115 6116 3149
rect 6050 3081 6116 3115
rect 6050 3047 6066 3081
rect 6100 3047 6116 3081
rect 6050 3038 6116 3047
rect 5651 2978 5705 2994
rect 5845 3013 6116 3038
rect 5845 3004 6066 3013
rect 5845 2990 5879 3004
rect 5651 2840 5685 2978
rect 5741 2956 5879 2990
rect 6050 2979 6066 3004
rect 6100 2979 6116 3013
rect 6156 3149 6206 3165
rect 6190 3115 6206 3149
rect 6250 3156 6266 3190
rect 6300 3156 6316 3190
rect 6250 3140 6316 3156
rect 6156 3106 6206 3115
rect 6354 3122 6420 3165
rect 6354 3106 6370 3122
rect 6156 3088 6370 3106
rect 6404 3088 6420 3122
rect 6156 3072 6420 3088
rect 6455 3125 6521 3263
rect 6455 3091 6471 3125
rect 6505 3091 6521 3125
rect 6455 3075 6521 3091
rect 6648 3149 6733 3165
rect 6648 3115 6664 3149
rect 6698 3115 6733 3149
rect 6156 3057 6206 3072
rect 6190 3023 6206 3057
rect 6648 3038 6733 3115
rect 6156 3007 6206 3023
rect 5947 2964 5993 2970
rect 5741 2940 5775 2956
rect 5719 2924 5775 2940
rect 5753 2890 5775 2924
rect 5947 2930 5953 2964
rect 5987 2930 5993 2964
rect 6050 2963 6116 2979
rect 6240 3004 6664 3038
rect 6698 3004 6733 3038
rect 6767 3149 6824 3165
rect 6767 3115 6783 3149
rect 6817 3115 6824 3149
rect 6767 3065 6824 3115
rect 6858 3151 6999 3263
rect 7185 3194 7251 3263
rect 7696 3259 7727 3293
rect 7761 3259 7823 3293
rect 7857 3259 7919 3293
rect 7953 3259 8015 3293
rect 8049 3259 8111 3293
rect 8145 3259 8207 3293
rect 8241 3259 8303 3293
rect 8337 3259 8399 3293
rect 8433 3259 8495 3293
rect 8529 3259 8591 3293
rect 8625 3259 8687 3293
rect 8721 3259 8783 3293
rect 8817 3259 8879 3293
rect 8913 3259 8975 3293
rect 9009 3259 9071 3293
rect 9105 3259 9167 3293
rect 9201 3259 9263 3293
rect 9297 3259 9359 3293
rect 9393 3259 9424 3293
rect 6858 3117 6874 3151
rect 6908 3117 6949 3151
rect 6983 3117 6999 3151
rect 6858 3114 6999 3117
rect 7034 3164 7098 3180
rect 7034 3130 7048 3164
rect 7082 3130 7098 3164
rect 7034 3065 7098 3130
rect 6767 3031 6783 3065
rect 6817 3054 7098 3065
rect 6817 3031 7048 3054
rect 7032 3020 7048 3031
rect 7082 3020 7098 3054
rect 7032 3004 7098 3020
rect 7185 3160 7201 3194
rect 7235 3160 7251 3194
rect 7185 3111 7251 3160
rect 7185 3077 7201 3111
rect 7235 3077 7251 3111
rect 7185 3028 7251 3077
rect 6240 2973 6274 3004
rect 5947 2929 5993 2930
rect 6150 2939 6274 2973
rect 6699 2997 6733 3004
rect 6402 2964 6473 2970
rect 6150 2929 6184 2939
rect 5719 2874 5775 2890
rect 5651 2824 5707 2840
rect 5651 2790 5673 2824
rect 5651 2734 5707 2790
rect 5651 2700 5673 2734
rect 5741 2764 5775 2874
rect 5811 2908 5877 2922
rect 5811 2874 5827 2908
rect 5861 2874 5877 2908
rect 5811 2858 5877 2874
rect 5947 2913 6057 2929
rect 5947 2879 6007 2913
rect 6041 2879 6057 2913
rect 5947 2866 6057 2879
rect 6099 2913 6184 2929
rect 6099 2879 6115 2913
rect 6149 2879 6184 2913
rect 6402 2930 6433 2964
rect 6467 2930 6473 2964
rect 6402 2913 6473 2930
rect 6099 2866 6184 2879
rect 6294 2889 6360 2905
rect 5843 2832 5877 2858
rect 6294 2855 6310 2889
rect 6344 2855 6360 2889
rect 6402 2879 6418 2913
rect 6452 2879 6473 2913
rect 6619 2964 6665 2970
rect 6619 2930 6625 2964
rect 6659 2930 6665 2964
rect 6699 2963 6944 2997
rect 7185 2994 7201 3028
rect 7235 2994 7251 3028
rect 7185 2978 7251 2994
rect 7291 3194 7342 3210
rect 7325 3160 7342 3194
rect 7291 3111 7342 3160
rect 7325 3077 7342 3111
rect 7291 3028 7342 3077
rect 7325 2994 7342 3028
rect 6619 2929 6665 2930
rect 6619 2913 6762 2929
rect 6402 2866 6473 2879
rect 6510 2890 6576 2905
rect 6510 2889 6532 2890
rect 6294 2832 6360 2855
rect 6510 2855 6526 2889
rect 6566 2856 6576 2890
rect 6619 2879 6712 2913
rect 6746 2879 6762 2913
rect 6619 2869 6762 2879
rect 6796 2913 6876 2929
rect 6796 2879 6826 2913
rect 6860 2879 6876 2913
rect 6796 2878 6876 2879
rect 6560 2855 6576 2856
rect 6510 2835 6576 2855
rect 6796 2835 6830 2878
rect 6910 2844 6944 2963
rect 6994 2934 7128 2970
rect 6994 2928 7056 2934
rect 7096 2928 7128 2934
rect 6994 2894 7010 2928
rect 7044 2894 7056 2928
rect 7112 2894 7128 2928
rect 7291 2954 7342 2994
rect 7713 3190 7767 3206
rect 7713 3156 7733 3190
rect 7713 3107 7767 3156
rect 7713 3073 7733 3107
rect 7713 3024 7767 3073
rect 7713 2990 7733 3024
rect 7807 3190 7873 3259
rect 7807 3156 7823 3190
rect 7857 3156 7873 3190
rect 8312 3186 8378 3259
rect 7807 3122 7873 3156
rect 7807 3088 7823 3122
rect 7857 3088 7873 3122
rect 7807 3054 7873 3088
rect 7807 3020 7823 3054
rect 7857 3020 7873 3054
rect 8112 3145 8178 3161
rect 8112 3111 8128 3145
rect 8162 3111 8178 3145
rect 8112 3077 8178 3111
rect 8112 3043 8128 3077
rect 8162 3043 8178 3077
rect 8112 3034 8178 3043
rect 7713 2974 7767 2990
rect 7907 3009 8178 3034
rect 7907 3000 8128 3009
rect 7907 2986 7941 3000
rect 6994 2892 7056 2894
rect 7096 2892 7128 2894
rect 6994 2878 7128 2892
rect 7176 2908 7242 2924
rect 7176 2874 7192 2908
rect 7226 2874 7242 2908
rect 7176 2844 7242 2874
rect 6510 2832 6830 2835
rect 5843 2801 6830 2832
rect 6864 2810 7242 2844
rect 7291 2920 7310 2954
rect 7291 2840 7342 2920
rect 7276 2824 7342 2840
rect 5843 2798 6576 2801
rect 6864 2767 6898 2810
rect 7276 2790 7292 2824
rect 7326 2790 7342 2824
rect 5741 2741 6088 2764
rect 5741 2730 6038 2741
rect 5651 2684 5707 2700
rect 6022 2707 6038 2730
rect 6072 2707 6088 2741
rect 5759 2662 5777 2696
rect 5811 2662 5830 2696
rect 6022 2685 6088 2707
rect 6130 2748 6416 2764
rect 6130 2714 6154 2748
rect 6188 2730 6366 2748
rect 6188 2714 6212 2730
rect 6130 2698 6212 2714
rect 6350 2714 6366 2730
rect 6400 2714 6416 2748
rect 6350 2698 6416 2714
rect 6450 2740 6545 2756
rect 6450 2706 6480 2740
rect 6514 2706 6545 2740
rect 3560 2599 3591 2633
rect 3625 2599 3687 2633
rect 3721 2599 3783 2633
rect 3817 2599 3879 2633
rect 3913 2599 3975 2633
rect 4009 2599 4071 2633
rect 4105 2599 4167 2633
rect 4201 2599 4263 2633
rect 4297 2599 4359 2633
rect 4393 2599 4455 2633
rect 4489 2599 4551 2633
rect 4585 2599 4647 2633
rect 4681 2599 4743 2633
rect 4777 2599 4839 2633
rect 4873 2599 4935 2633
rect 4969 2599 5031 2633
rect 5065 2599 5127 2633
rect 5161 2599 5223 2633
rect 5257 2599 5288 2633
rect 5759 2631 5830 2662
rect 6248 2662 6264 2696
rect 6298 2662 6314 2696
rect 6248 2631 6314 2662
rect 6450 2631 6545 2706
rect 6643 2751 6898 2767
rect 6643 2717 6659 2751
rect 6693 2733 6898 2751
rect 6932 2760 7152 2776
rect 6932 2742 7102 2760
rect 6693 2717 6709 2733
rect 6643 2701 6709 2717
rect 6932 2699 6966 2742
rect 7086 2726 7102 2742
rect 7136 2726 7152 2760
rect 7086 2710 7152 2726
rect 7190 2752 7240 2768
rect 7190 2718 7206 2752
rect 6745 2665 6761 2699
rect 6795 2665 6855 2699
rect 6889 2665 6966 2699
rect 7000 2692 7050 2708
rect 7034 2658 7050 2692
rect 7000 2631 7050 2658
rect 7190 2631 7240 2718
rect 7276 2734 7342 2790
rect 7276 2700 7292 2734
rect 7326 2700 7342 2734
rect 7276 2684 7342 2700
rect 7713 2836 7747 2974
rect 7803 2952 7941 2986
rect 8112 2975 8128 3000
rect 8162 2975 8178 3009
rect 8218 3145 8268 3161
rect 8252 3111 8268 3145
rect 8312 3152 8328 3186
rect 8362 3152 8378 3186
rect 8312 3136 8378 3152
rect 8218 3102 8268 3111
rect 8416 3118 8482 3161
rect 8416 3102 8432 3118
rect 8218 3084 8432 3102
rect 8466 3084 8482 3118
rect 8218 3068 8482 3084
rect 8517 3121 8583 3259
rect 8517 3087 8533 3121
rect 8567 3087 8583 3121
rect 8517 3071 8583 3087
rect 8710 3145 8795 3161
rect 8710 3111 8726 3145
rect 8760 3111 8795 3145
rect 8218 3053 8268 3068
rect 8252 3019 8268 3053
rect 8710 3034 8795 3111
rect 8218 3003 8268 3019
rect 8009 2960 8055 2966
rect 7803 2936 7837 2952
rect 7781 2920 7837 2936
rect 7815 2886 7837 2920
rect 8009 2926 8015 2960
rect 8049 2926 8055 2960
rect 8112 2959 8178 2975
rect 8302 3000 8726 3034
rect 8760 3000 8795 3034
rect 8829 3145 8886 3161
rect 8829 3111 8845 3145
rect 8879 3111 8886 3145
rect 8829 3061 8886 3111
rect 8920 3147 9061 3259
rect 9247 3190 9313 3259
rect 9756 3255 9787 3289
rect 9821 3255 9883 3289
rect 9917 3255 9979 3289
rect 10013 3255 10075 3289
rect 10109 3255 10171 3289
rect 10205 3255 10267 3289
rect 10301 3255 10363 3289
rect 10397 3255 10459 3289
rect 10493 3255 10555 3289
rect 10589 3255 10651 3289
rect 10685 3255 10747 3289
rect 10781 3255 10843 3289
rect 10877 3255 10939 3289
rect 10973 3255 11035 3289
rect 11069 3255 11131 3289
rect 11165 3255 11227 3289
rect 11261 3255 11323 3289
rect 11357 3255 11419 3289
rect 11453 3255 11484 3289
rect 8920 3113 8936 3147
rect 8970 3113 9011 3147
rect 9045 3113 9061 3147
rect 8920 3110 9061 3113
rect 9096 3160 9160 3176
rect 9096 3126 9110 3160
rect 9144 3126 9160 3160
rect 9096 3061 9160 3126
rect 8829 3027 8845 3061
rect 8879 3050 9160 3061
rect 8879 3027 9110 3050
rect 9094 3016 9110 3027
rect 9144 3016 9160 3050
rect 9094 3000 9160 3016
rect 9247 3156 9263 3190
rect 9297 3156 9313 3190
rect 9247 3107 9313 3156
rect 9247 3073 9263 3107
rect 9297 3073 9313 3107
rect 9247 3024 9313 3073
rect 8302 2969 8336 3000
rect 8009 2925 8055 2926
rect 8212 2935 8336 2969
rect 8761 2993 8795 3000
rect 8464 2960 8535 2966
rect 8212 2925 8246 2935
rect 7781 2870 7837 2886
rect 7713 2820 7769 2836
rect 7713 2786 7735 2820
rect 7713 2730 7769 2786
rect 7713 2696 7735 2730
rect 7803 2760 7837 2870
rect 7873 2904 7939 2918
rect 7873 2870 7889 2904
rect 7923 2870 7939 2904
rect 7873 2854 7939 2870
rect 8009 2909 8119 2925
rect 8009 2875 8069 2909
rect 8103 2875 8119 2909
rect 8009 2862 8119 2875
rect 8161 2909 8246 2925
rect 8161 2875 8177 2909
rect 8211 2875 8246 2909
rect 8464 2926 8495 2960
rect 8529 2926 8535 2960
rect 8464 2909 8535 2926
rect 8161 2862 8246 2875
rect 8356 2885 8422 2901
rect 7905 2828 7939 2854
rect 8356 2851 8372 2885
rect 8406 2851 8422 2885
rect 8464 2875 8480 2909
rect 8514 2875 8535 2909
rect 8681 2960 8727 2966
rect 8681 2926 8687 2960
rect 8721 2926 8727 2960
rect 8761 2959 9006 2993
rect 9247 2990 9263 3024
rect 9297 2990 9313 3024
rect 9247 2974 9313 2990
rect 9353 3190 9404 3206
rect 9387 3156 9404 3190
rect 9353 3107 9404 3156
rect 9387 3073 9404 3107
rect 9353 3024 9404 3073
rect 9387 2990 9404 3024
rect 8681 2925 8727 2926
rect 8681 2909 8824 2925
rect 8464 2862 8535 2875
rect 8572 2886 8638 2901
rect 8572 2885 8594 2886
rect 8356 2828 8422 2851
rect 8572 2851 8588 2885
rect 8628 2852 8638 2886
rect 8681 2875 8774 2909
rect 8808 2875 8824 2909
rect 8681 2865 8824 2875
rect 8858 2909 8938 2925
rect 8858 2875 8888 2909
rect 8922 2875 8938 2909
rect 8858 2874 8938 2875
rect 8622 2851 8638 2852
rect 8572 2831 8638 2851
rect 8858 2831 8892 2874
rect 8972 2840 9006 2959
rect 9056 2930 9190 2966
rect 9056 2924 9118 2930
rect 9158 2924 9190 2930
rect 9056 2890 9072 2924
rect 9106 2890 9118 2924
rect 9174 2890 9190 2924
rect 9353 2944 9404 2990
rect 9056 2888 9118 2890
rect 9158 2888 9190 2890
rect 9056 2874 9190 2888
rect 9238 2904 9304 2920
rect 9238 2870 9254 2904
rect 9288 2870 9304 2904
rect 9238 2840 9304 2870
rect 8572 2828 8892 2831
rect 7905 2797 8892 2828
rect 8926 2806 9304 2840
rect 9353 2910 9366 2944
rect 9402 2910 9404 2944
rect 9353 2836 9404 2910
rect 9338 2820 9404 2836
rect 7905 2794 8638 2797
rect 8926 2763 8960 2806
rect 9338 2786 9354 2820
rect 9388 2786 9404 2820
rect 7803 2737 8150 2760
rect 7803 2726 8100 2737
rect 7713 2680 7769 2696
rect 8084 2703 8100 2726
rect 8134 2703 8150 2737
rect 7821 2658 7839 2692
rect 7873 2658 7892 2692
rect 8084 2681 8150 2703
rect 8192 2744 8478 2760
rect 8192 2710 8216 2744
rect 8250 2726 8428 2744
rect 8250 2710 8274 2726
rect 8192 2694 8274 2710
rect 8412 2710 8428 2726
rect 8462 2710 8478 2744
rect 8412 2694 8478 2710
rect 8512 2736 8607 2752
rect 8512 2702 8542 2736
rect 8576 2702 8607 2736
rect 5634 2597 5665 2631
rect 5699 2597 5761 2631
rect 5795 2597 5857 2631
rect 5891 2597 5953 2631
rect 5987 2597 6049 2631
rect 6083 2597 6145 2631
rect 6179 2597 6241 2631
rect 6275 2597 6337 2631
rect 6371 2597 6433 2631
rect 6467 2597 6529 2631
rect 6563 2597 6625 2631
rect 6659 2597 6721 2631
rect 6755 2597 6817 2631
rect 6851 2597 6913 2631
rect 6947 2597 7009 2631
rect 7043 2597 7105 2631
rect 7139 2597 7201 2631
rect 7235 2597 7297 2631
rect 7331 2597 7362 2631
rect 7821 2627 7892 2658
rect 8310 2658 8326 2692
rect 8360 2658 8376 2692
rect 8310 2627 8376 2658
rect 8512 2627 8607 2702
rect 8705 2747 8960 2763
rect 8705 2713 8721 2747
rect 8755 2729 8960 2747
rect 8994 2756 9214 2772
rect 8994 2738 9164 2756
rect 8755 2713 8771 2729
rect 8705 2697 8771 2713
rect 8994 2695 9028 2738
rect 9148 2722 9164 2738
rect 9198 2722 9214 2756
rect 9148 2706 9214 2722
rect 9252 2748 9302 2764
rect 9252 2714 9268 2748
rect 8807 2661 8823 2695
rect 8857 2661 8917 2695
rect 8951 2661 9028 2695
rect 9062 2688 9112 2704
rect 9096 2654 9112 2688
rect 9062 2627 9112 2654
rect 9252 2627 9302 2714
rect 9338 2730 9404 2786
rect 9338 2696 9354 2730
rect 9388 2696 9404 2730
rect 9338 2680 9404 2696
rect 9773 3186 9827 3202
rect 9773 3152 9793 3186
rect 9773 3103 9827 3152
rect 9773 3069 9793 3103
rect 9773 3020 9827 3069
rect 9773 2986 9793 3020
rect 9867 3186 9933 3255
rect 9867 3152 9883 3186
rect 9917 3152 9933 3186
rect 10372 3182 10438 3255
rect 9867 3118 9933 3152
rect 9867 3084 9883 3118
rect 9917 3084 9933 3118
rect 9867 3050 9933 3084
rect 9867 3016 9883 3050
rect 9917 3016 9933 3050
rect 10172 3141 10238 3157
rect 10172 3107 10188 3141
rect 10222 3107 10238 3141
rect 10172 3073 10238 3107
rect 10172 3039 10188 3073
rect 10222 3039 10238 3073
rect 10172 3030 10238 3039
rect 9773 2970 9827 2986
rect 9967 3005 10238 3030
rect 9967 2996 10188 3005
rect 9967 2982 10001 2996
rect 9773 2832 9807 2970
rect 9863 2948 10001 2982
rect 10172 2971 10188 2996
rect 10222 2971 10238 3005
rect 10278 3141 10328 3157
rect 10312 3107 10328 3141
rect 10372 3148 10388 3182
rect 10422 3148 10438 3182
rect 10372 3132 10438 3148
rect 10278 3098 10328 3107
rect 10476 3114 10542 3157
rect 10476 3098 10492 3114
rect 10278 3080 10492 3098
rect 10526 3080 10542 3114
rect 10278 3064 10542 3080
rect 10577 3117 10643 3255
rect 10577 3083 10593 3117
rect 10627 3083 10643 3117
rect 10577 3067 10643 3083
rect 10770 3141 10855 3157
rect 10770 3107 10786 3141
rect 10820 3107 10855 3141
rect 10278 3049 10328 3064
rect 10312 3015 10328 3049
rect 10770 3030 10855 3107
rect 10278 2999 10328 3015
rect 10069 2956 10115 2962
rect 9863 2932 9897 2948
rect 9841 2916 9897 2932
rect 9875 2882 9897 2916
rect 10069 2922 10075 2956
rect 10109 2922 10115 2956
rect 10172 2955 10238 2971
rect 10362 2996 10786 3030
rect 10820 2996 10855 3030
rect 10889 3141 10946 3157
rect 10889 3107 10905 3141
rect 10939 3107 10946 3141
rect 10889 3057 10946 3107
rect 10980 3143 11121 3255
rect 11307 3186 11373 3255
rect 11818 3251 11849 3285
rect 11883 3251 11945 3285
rect 11979 3251 12041 3285
rect 12075 3251 12137 3285
rect 12171 3251 12233 3285
rect 12267 3251 12329 3285
rect 12363 3251 12425 3285
rect 12459 3251 12521 3285
rect 12555 3251 12617 3285
rect 12651 3251 12713 3285
rect 12747 3251 12809 3285
rect 12843 3251 12905 3285
rect 12939 3251 13001 3285
rect 13035 3251 13097 3285
rect 13131 3251 13193 3285
rect 13227 3251 13289 3285
rect 13323 3251 13385 3285
rect 13419 3251 13481 3285
rect 13515 3251 13546 3285
rect 10980 3109 10996 3143
rect 11030 3109 11071 3143
rect 11105 3109 11121 3143
rect 10980 3106 11121 3109
rect 11156 3156 11220 3172
rect 11156 3122 11170 3156
rect 11204 3122 11220 3156
rect 11156 3057 11220 3122
rect 10889 3023 10905 3057
rect 10939 3046 11220 3057
rect 10939 3023 11170 3046
rect 11154 3012 11170 3023
rect 11204 3012 11220 3046
rect 11154 2996 11220 3012
rect 11307 3152 11323 3186
rect 11357 3152 11373 3186
rect 11307 3103 11373 3152
rect 11307 3069 11323 3103
rect 11357 3069 11373 3103
rect 11307 3020 11373 3069
rect 10362 2965 10396 2996
rect 10069 2921 10115 2922
rect 10272 2931 10396 2965
rect 10821 2989 10855 2996
rect 10524 2956 10595 2962
rect 10272 2921 10306 2931
rect 9841 2866 9897 2882
rect 9773 2816 9829 2832
rect 9773 2782 9795 2816
rect 9773 2726 9829 2782
rect 9773 2692 9795 2726
rect 9863 2756 9897 2866
rect 9933 2900 9999 2914
rect 9933 2866 9949 2900
rect 9983 2866 9999 2900
rect 9933 2850 9999 2866
rect 10069 2905 10179 2921
rect 10069 2871 10129 2905
rect 10163 2871 10179 2905
rect 10069 2858 10179 2871
rect 10221 2905 10306 2921
rect 10221 2871 10237 2905
rect 10271 2871 10306 2905
rect 10524 2922 10555 2956
rect 10589 2922 10595 2956
rect 10524 2905 10595 2922
rect 10221 2858 10306 2871
rect 10416 2881 10482 2897
rect 9965 2824 9999 2850
rect 10416 2847 10432 2881
rect 10466 2847 10482 2881
rect 10524 2871 10540 2905
rect 10574 2871 10595 2905
rect 10741 2956 10787 2962
rect 10741 2922 10747 2956
rect 10781 2922 10787 2956
rect 10821 2955 11066 2989
rect 11307 2986 11323 3020
rect 11357 2986 11373 3020
rect 11307 2970 11373 2986
rect 11413 3186 11464 3202
rect 11447 3152 11464 3186
rect 11413 3103 11464 3152
rect 11447 3069 11464 3103
rect 11413 3020 11464 3069
rect 11447 2986 11464 3020
rect 10741 2921 10787 2922
rect 10741 2905 10884 2921
rect 10524 2858 10595 2871
rect 10632 2882 10698 2897
rect 10632 2881 10654 2882
rect 10416 2824 10482 2847
rect 10632 2847 10648 2881
rect 10688 2848 10698 2882
rect 10741 2871 10834 2905
rect 10868 2871 10884 2905
rect 10741 2861 10884 2871
rect 10918 2905 10998 2921
rect 10918 2871 10948 2905
rect 10982 2871 10998 2905
rect 10918 2870 10998 2871
rect 10682 2847 10698 2848
rect 10632 2827 10698 2847
rect 10918 2827 10952 2870
rect 11032 2836 11066 2955
rect 11116 2926 11250 2962
rect 11116 2920 11178 2926
rect 11218 2920 11250 2926
rect 11116 2886 11132 2920
rect 11166 2886 11178 2920
rect 11234 2886 11250 2920
rect 11413 2946 11464 2986
rect 11835 3182 11889 3198
rect 11835 3148 11855 3182
rect 11835 3099 11889 3148
rect 11835 3065 11855 3099
rect 11835 3016 11889 3065
rect 11835 2982 11855 3016
rect 11929 3182 11995 3251
rect 11929 3148 11945 3182
rect 11979 3148 11995 3182
rect 12434 3178 12500 3251
rect 11929 3114 11995 3148
rect 11929 3080 11945 3114
rect 11979 3080 11995 3114
rect 11929 3046 11995 3080
rect 11929 3012 11945 3046
rect 11979 3012 11995 3046
rect 12234 3137 12300 3153
rect 12234 3103 12250 3137
rect 12284 3103 12300 3137
rect 12234 3069 12300 3103
rect 12234 3035 12250 3069
rect 12284 3035 12300 3069
rect 12234 3026 12300 3035
rect 11835 2966 11889 2982
rect 12029 3001 12300 3026
rect 12029 2992 12250 3001
rect 12029 2978 12063 2992
rect 11116 2884 11178 2886
rect 11218 2884 11250 2886
rect 11116 2870 11250 2884
rect 11298 2900 11364 2916
rect 11298 2866 11314 2900
rect 11348 2866 11364 2900
rect 11298 2836 11364 2866
rect 10632 2824 10952 2827
rect 9965 2793 10952 2824
rect 10986 2802 11364 2836
rect 11413 2912 11432 2946
rect 11413 2832 11464 2912
rect 11398 2816 11464 2832
rect 9965 2790 10698 2793
rect 10986 2759 11020 2802
rect 11398 2782 11414 2816
rect 11448 2782 11464 2816
rect 9863 2733 10210 2756
rect 9863 2722 10160 2733
rect 9773 2676 9829 2692
rect 10144 2699 10160 2722
rect 10194 2699 10210 2733
rect 9881 2654 9899 2688
rect 9933 2654 9952 2688
rect 10144 2677 10210 2699
rect 10252 2740 10538 2756
rect 10252 2706 10276 2740
rect 10310 2722 10488 2740
rect 10310 2706 10334 2722
rect 10252 2690 10334 2706
rect 10472 2706 10488 2722
rect 10522 2706 10538 2740
rect 10472 2690 10538 2706
rect 10572 2732 10667 2748
rect 10572 2698 10602 2732
rect 10636 2698 10667 2732
rect 7696 2593 7727 2627
rect 7761 2593 7823 2627
rect 7857 2593 7919 2627
rect 7953 2593 8015 2627
rect 8049 2593 8111 2627
rect 8145 2593 8207 2627
rect 8241 2593 8303 2627
rect 8337 2593 8399 2627
rect 8433 2593 8495 2627
rect 8529 2593 8591 2627
rect 8625 2593 8687 2627
rect 8721 2593 8783 2627
rect 8817 2593 8879 2627
rect 8913 2593 8975 2627
rect 9009 2593 9071 2627
rect 9105 2593 9167 2627
rect 9201 2593 9263 2627
rect 9297 2593 9359 2627
rect 9393 2593 9424 2627
rect 9881 2623 9952 2654
rect 10370 2654 10386 2688
rect 10420 2654 10436 2688
rect 10370 2623 10436 2654
rect 10572 2623 10667 2698
rect 10765 2743 11020 2759
rect 10765 2709 10781 2743
rect 10815 2725 11020 2743
rect 11054 2752 11274 2768
rect 11054 2734 11224 2752
rect 10815 2709 10831 2725
rect 10765 2693 10831 2709
rect 11054 2691 11088 2734
rect 11208 2718 11224 2734
rect 11258 2718 11274 2752
rect 11208 2702 11274 2718
rect 11312 2744 11362 2760
rect 11312 2710 11328 2744
rect 10867 2657 10883 2691
rect 10917 2657 10977 2691
rect 11011 2657 11088 2691
rect 11122 2684 11172 2700
rect 11156 2650 11172 2684
rect 11122 2623 11172 2650
rect 11312 2623 11362 2710
rect 11398 2726 11464 2782
rect 11398 2692 11414 2726
rect 11448 2692 11464 2726
rect 11398 2676 11464 2692
rect 11835 2828 11869 2966
rect 11925 2944 12063 2978
rect 12234 2967 12250 2992
rect 12284 2967 12300 3001
rect 12340 3137 12390 3153
rect 12374 3103 12390 3137
rect 12434 3144 12450 3178
rect 12484 3144 12500 3178
rect 12434 3128 12500 3144
rect 12340 3094 12390 3103
rect 12538 3110 12604 3153
rect 12538 3094 12554 3110
rect 12340 3076 12554 3094
rect 12588 3076 12604 3110
rect 12340 3060 12604 3076
rect 12639 3113 12705 3251
rect 12639 3079 12655 3113
rect 12689 3079 12705 3113
rect 12639 3063 12705 3079
rect 12832 3137 12917 3153
rect 12832 3103 12848 3137
rect 12882 3103 12917 3137
rect 12340 3045 12390 3060
rect 12374 3011 12390 3045
rect 12832 3026 12917 3103
rect 12340 2995 12390 3011
rect 12131 2952 12177 2958
rect 11925 2928 11959 2944
rect 11903 2912 11959 2928
rect 11937 2878 11959 2912
rect 12131 2918 12137 2952
rect 12171 2918 12177 2952
rect 12234 2951 12300 2967
rect 12424 2992 12848 3026
rect 12882 2992 12917 3026
rect 12951 3137 13008 3153
rect 12951 3103 12967 3137
rect 13001 3103 13008 3137
rect 12951 3053 13008 3103
rect 13042 3139 13183 3251
rect 13369 3182 13435 3251
rect 13892 3249 13923 3283
rect 13957 3249 14019 3283
rect 14053 3249 14115 3283
rect 14149 3249 14211 3283
rect 14245 3249 14307 3283
rect 14341 3249 14403 3283
rect 14437 3249 14499 3283
rect 14533 3249 14595 3283
rect 14629 3249 14691 3283
rect 14725 3249 14787 3283
rect 14821 3249 14883 3283
rect 14917 3249 14979 3283
rect 15013 3249 15075 3283
rect 15109 3249 15171 3283
rect 15205 3249 15267 3283
rect 15301 3249 15363 3283
rect 15397 3249 15459 3283
rect 15493 3249 15555 3283
rect 15589 3249 15620 3283
rect 13042 3105 13058 3139
rect 13092 3105 13133 3139
rect 13167 3105 13183 3139
rect 13042 3102 13183 3105
rect 13218 3152 13282 3168
rect 13218 3118 13232 3152
rect 13266 3118 13282 3152
rect 13218 3053 13282 3118
rect 12951 3019 12967 3053
rect 13001 3042 13282 3053
rect 13001 3019 13232 3042
rect 13216 3008 13232 3019
rect 13266 3008 13282 3042
rect 13216 2992 13282 3008
rect 13369 3148 13385 3182
rect 13419 3148 13435 3182
rect 13369 3099 13435 3148
rect 13369 3065 13385 3099
rect 13419 3065 13435 3099
rect 13369 3016 13435 3065
rect 12424 2961 12458 2992
rect 12131 2917 12177 2918
rect 12334 2927 12458 2961
rect 12883 2985 12917 2992
rect 12586 2952 12657 2958
rect 12334 2917 12368 2927
rect 11903 2862 11959 2878
rect 11835 2812 11891 2828
rect 11835 2778 11857 2812
rect 11835 2722 11891 2778
rect 11835 2688 11857 2722
rect 11925 2752 11959 2862
rect 11995 2896 12061 2910
rect 11995 2862 12011 2896
rect 12045 2862 12061 2896
rect 11995 2846 12061 2862
rect 12131 2901 12241 2917
rect 12131 2867 12191 2901
rect 12225 2867 12241 2901
rect 12131 2854 12241 2867
rect 12283 2901 12368 2917
rect 12283 2867 12299 2901
rect 12333 2867 12368 2901
rect 12586 2918 12617 2952
rect 12651 2918 12657 2952
rect 12586 2901 12657 2918
rect 12283 2854 12368 2867
rect 12478 2877 12544 2893
rect 12027 2820 12061 2846
rect 12478 2843 12494 2877
rect 12528 2843 12544 2877
rect 12586 2867 12602 2901
rect 12636 2867 12657 2901
rect 12803 2952 12849 2958
rect 12803 2918 12809 2952
rect 12843 2918 12849 2952
rect 12883 2951 13128 2985
rect 13369 2982 13385 3016
rect 13419 2982 13435 3016
rect 13369 2966 13435 2982
rect 13475 3182 13526 3198
rect 13509 3148 13526 3182
rect 13475 3099 13526 3148
rect 13509 3065 13526 3099
rect 13475 3016 13526 3065
rect 13509 2982 13526 3016
rect 12803 2917 12849 2918
rect 12803 2901 12946 2917
rect 12586 2854 12657 2867
rect 12694 2878 12760 2893
rect 12694 2877 12716 2878
rect 12478 2820 12544 2843
rect 12694 2843 12710 2877
rect 12750 2844 12760 2878
rect 12803 2867 12896 2901
rect 12930 2867 12946 2901
rect 12803 2857 12946 2867
rect 12980 2901 13060 2917
rect 12980 2867 13010 2901
rect 13044 2867 13060 2901
rect 12980 2866 13060 2867
rect 12744 2843 12760 2844
rect 12694 2823 12760 2843
rect 12980 2823 13014 2866
rect 13094 2832 13128 2951
rect 13178 2922 13312 2958
rect 13178 2916 13240 2922
rect 13280 2916 13312 2922
rect 13178 2882 13194 2916
rect 13228 2882 13240 2916
rect 13296 2882 13312 2916
rect 13475 2948 13526 2982
rect 13475 2914 13490 2948
rect 13178 2880 13240 2882
rect 13280 2880 13312 2882
rect 13178 2866 13312 2880
rect 13360 2896 13426 2912
rect 13360 2862 13376 2896
rect 13410 2862 13426 2896
rect 13360 2832 13426 2862
rect 12694 2820 13014 2823
rect 12027 2789 13014 2820
rect 13048 2798 13426 2832
rect 13475 2828 13526 2914
rect 13460 2812 13526 2828
rect 12027 2786 12760 2789
rect 13048 2755 13082 2798
rect 13460 2778 13476 2812
rect 13510 2778 13526 2812
rect 11925 2729 12272 2752
rect 11925 2718 12222 2729
rect 11835 2672 11891 2688
rect 12206 2695 12222 2718
rect 12256 2695 12272 2729
rect 11943 2650 11961 2684
rect 11995 2650 12014 2684
rect 12206 2673 12272 2695
rect 12314 2736 12600 2752
rect 12314 2702 12338 2736
rect 12372 2718 12550 2736
rect 12372 2702 12396 2718
rect 12314 2686 12396 2702
rect 12534 2702 12550 2718
rect 12584 2702 12600 2736
rect 12534 2686 12600 2702
rect 12634 2728 12729 2744
rect 12634 2694 12664 2728
rect 12698 2694 12729 2728
rect 9756 2589 9787 2623
rect 9821 2589 9883 2623
rect 9917 2589 9979 2623
rect 10013 2589 10075 2623
rect 10109 2589 10171 2623
rect 10205 2589 10267 2623
rect 10301 2589 10363 2623
rect 10397 2589 10459 2623
rect 10493 2589 10555 2623
rect 10589 2589 10651 2623
rect 10685 2589 10747 2623
rect 10781 2589 10843 2623
rect 10877 2589 10939 2623
rect 10973 2589 11035 2623
rect 11069 2589 11131 2623
rect 11165 2589 11227 2623
rect 11261 2589 11323 2623
rect 11357 2589 11419 2623
rect 11453 2589 11484 2623
rect 11943 2619 12014 2650
rect 12432 2650 12448 2684
rect 12482 2650 12498 2684
rect 12432 2619 12498 2650
rect 12634 2619 12729 2694
rect 12827 2739 13082 2755
rect 12827 2705 12843 2739
rect 12877 2721 13082 2739
rect 13116 2748 13336 2764
rect 13116 2730 13286 2748
rect 12877 2705 12893 2721
rect 12827 2689 12893 2705
rect 13116 2687 13150 2730
rect 13270 2714 13286 2730
rect 13320 2714 13336 2748
rect 13270 2698 13336 2714
rect 13374 2740 13424 2756
rect 13374 2706 13390 2740
rect 12929 2653 12945 2687
rect 12979 2653 13039 2687
rect 13073 2653 13150 2687
rect 13184 2680 13234 2696
rect 13218 2646 13234 2680
rect 13184 2619 13234 2646
rect 13374 2619 13424 2706
rect 13460 2722 13526 2778
rect 13460 2688 13476 2722
rect 13510 2688 13526 2722
rect 13460 2672 13526 2688
rect 13909 3180 13963 3196
rect 13909 3146 13929 3180
rect 13909 3097 13963 3146
rect 13909 3063 13929 3097
rect 13909 3014 13963 3063
rect 13909 2980 13929 3014
rect 14003 3180 14069 3249
rect 14003 3146 14019 3180
rect 14053 3146 14069 3180
rect 14508 3176 14574 3249
rect 14003 3112 14069 3146
rect 14003 3078 14019 3112
rect 14053 3078 14069 3112
rect 14003 3044 14069 3078
rect 14003 3010 14019 3044
rect 14053 3010 14069 3044
rect 14308 3135 14374 3151
rect 14308 3101 14324 3135
rect 14358 3101 14374 3135
rect 14308 3067 14374 3101
rect 14308 3033 14324 3067
rect 14358 3033 14374 3067
rect 14308 3024 14374 3033
rect 13909 2964 13963 2980
rect 14103 2999 14374 3024
rect 14103 2990 14324 2999
rect 14103 2976 14137 2990
rect 13909 2826 13943 2964
rect 13999 2942 14137 2976
rect 14308 2965 14324 2990
rect 14358 2965 14374 2999
rect 14414 3135 14464 3151
rect 14448 3101 14464 3135
rect 14508 3142 14524 3176
rect 14558 3142 14574 3176
rect 14508 3126 14574 3142
rect 14414 3092 14464 3101
rect 14612 3108 14678 3151
rect 14612 3092 14628 3108
rect 14414 3074 14628 3092
rect 14662 3074 14678 3108
rect 14414 3058 14678 3074
rect 14713 3111 14779 3249
rect 14713 3077 14729 3111
rect 14763 3077 14779 3111
rect 14713 3061 14779 3077
rect 14906 3135 14991 3151
rect 14906 3101 14922 3135
rect 14956 3101 14991 3135
rect 14414 3043 14464 3058
rect 14448 3009 14464 3043
rect 14906 3024 14991 3101
rect 14414 2993 14464 3009
rect 14205 2950 14251 2956
rect 13999 2926 14033 2942
rect 13977 2910 14033 2926
rect 14011 2876 14033 2910
rect 14205 2916 14211 2950
rect 14245 2916 14251 2950
rect 14308 2949 14374 2965
rect 14498 2990 14922 3024
rect 14956 2990 14991 3024
rect 15025 3135 15082 3151
rect 15025 3101 15041 3135
rect 15075 3101 15082 3135
rect 15025 3051 15082 3101
rect 15116 3137 15257 3249
rect 15443 3180 15509 3249
rect 15954 3245 15985 3279
rect 16019 3245 16081 3279
rect 16115 3245 16177 3279
rect 16211 3245 16273 3279
rect 16307 3245 16369 3279
rect 16403 3245 16465 3279
rect 16499 3245 16561 3279
rect 16595 3245 16657 3279
rect 16691 3245 16753 3279
rect 16787 3245 16849 3279
rect 16883 3245 16945 3279
rect 16979 3245 17041 3279
rect 17075 3245 17137 3279
rect 17171 3245 17233 3279
rect 17267 3245 17329 3279
rect 17363 3245 17425 3279
rect 17459 3245 17521 3279
rect 17555 3245 17617 3279
rect 17651 3245 17682 3279
rect 15116 3103 15132 3137
rect 15166 3103 15207 3137
rect 15241 3103 15257 3137
rect 15116 3100 15257 3103
rect 15292 3150 15356 3166
rect 15292 3116 15306 3150
rect 15340 3116 15356 3150
rect 15292 3051 15356 3116
rect 15025 3017 15041 3051
rect 15075 3040 15356 3051
rect 15075 3017 15306 3040
rect 15290 3006 15306 3017
rect 15340 3006 15356 3040
rect 15290 2990 15356 3006
rect 15443 3146 15459 3180
rect 15493 3146 15509 3180
rect 15443 3097 15509 3146
rect 15443 3063 15459 3097
rect 15493 3063 15509 3097
rect 15443 3014 15509 3063
rect 14498 2959 14532 2990
rect 14205 2915 14251 2916
rect 14408 2925 14532 2959
rect 14957 2983 14991 2990
rect 14660 2950 14731 2956
rect 14408 2915 14442 2925
rect 13977 2860 14033 2876
rect 13909 2810 13965 2826
rect 13909 2776 13931 2810
rect 13909 2720 13965 2776
rect 13909 2686 13931 2720
rect 13999 2750 14033 2860
rect 14069 2894 14135 2908
rect 14069 2860 14085 2894
rect 14119 2860 14135 2894
rect 14069 2844 14135 2860
rect 14205 2899 14315 2915
rect 14205 2865 14265 2899
rect 14299 2865 14315 2899
rect 14205 2852 14315 2865
rect 14357 2899 14442 2915
rect 14357 2865 14373 2899
rect 14407 2865 14442 2899
rect 14660 2916 14691 2950
rect 14725 2916 14731 2950
rect 14660 2899 14731 2916
rect 14357 2852 14442 2865
rect 14552 2875 14618 2891
rect 14101 2818 14135 2844
rect 14552 2841 14568 2875
rect 14602 2841 14618 2875
rect 14660 2865 14676 2899
rect 14710 2865 14731 2899
rect 14877 2950 14923 2956
rect 14877 2916 14883 2950
rect 14917 2916 14923 2950
rect 14957 2949 15202 2983
rect 15443 2980 15459 3014
rect 15493 2980 15509 3014
rect 15443 2964 15509 2980
rect 15549 3180 15600 3196
rect 15583 3146 15600 3180
rect 15549 3097 15600 3146
rect 15583 3063 15600 3097
rect 15549 3014 15600 3063
rect 15583 2980 15600 3014
rect 14877 2915 14923 2916
rect 14877 2899 15020 2915
rect 14660 2852 14731 2865
rect 14768 2876 14834 2891
rect 14768 2875 14790 2876
rect 14552 2818 14618 2841
rect 14768 2841 14784 2875
rect 14824 2842 14834 2876
rect 14877 2865 14970 2899
rect 15004 2865 15020 2899
rect 14877 2855 15020 2865
rect 15054 2899 15134 2915
rect 15054 2865 15084 2899
rect 15118 2865 15134 2899
rect 15054 2864 15134 2865
rect 14818 2841 14834 2842
rect 14768 2821 14834 2841
rect 15054 2821 15088 2864
rect 15168 2830 15202 2949
rect 15252 2920 15386 2956
rect 15252 2914 15314 2920
rect 15354 2914 15386 2920
rect 15252 2880 15268 2914
rect 15302 2880 15314 2914
rect 15370 2880 15386 2914
rect 15549 2940 15600 2980
rect 15971 3176 16025 3192
rect 15971 3142 15991 3176
rect 15971 3093 16025 3142
rect 15971 3059 15991 3093
rect 15971 3010 16025 3059
rect 15971 2976 15991 3010
rect 16065 3176 16131 3245
rect 16065 3142 16081 3176
rect 16115 3142 16131 3176
rect 16570 3172 16636 3245
rect 16065 3108 16131 3142
rect 16065 3074 16081 3108
rect 16115 3074 16131 3108
rect 16065 3040 16131 3074
rect 16065 3006 16081 3040
rect 16115 3006 16131 3040
rect 16370 3131 16436 3147
rect 16370 3097 16386 3131
rect 16420 3097 16436 3131
rect 16370 3063 16436 3097
rect 16370 3029 16386 3063
rect 16420 3029 16436 3063
rect 16370 3020 16436 3029
rect 15971 2960 16025 2976
rect 16165 2995 16436 3020
rect 16165 2986 16386 2995
rect 16165 2972 16199 2986
rect 15252 2878 15314 2880
rect 15354 2878 15386 2880
rect 15252 2864 15386 2878
rect 15434 2894 15500 2910
rect 15434 2860 15450 2894
rect 15484 2860 15500 2894
rect 15434 2830 15500 2860
rect 14768 2818 15088 2821
rect 14101 2787 15088 2818
rect 15122 2796 15500 2830
rect 15549 2906 15568 2940
rect 15549 2826 15600 2906
rect 15534 2810 15600 2826
rect 14101 2784 14834 2787
rect 15122 2753 15156 2796
rect 15534 2776 15550 2810
rect 15584 2776 15600 2810
rect 13999 2727 14346 2750
rect 13999 2716 14296 2727
rect 13909 2670 13965 2686
rect 14280 2693 14296 2716
rect 14330 2693 14346 2727
rect 14017 2648 14035 2682
rect 14069 2648 14088 2682
rect 14280 2671 14346 2693
rect 14388 2734 14674 2750
rect 14388 2700 14412 2734
rect 14446 2716 14624 2734
rect 14446 2700 14470 2716
rect 14388 2684 14470 2700
rect 14608 2700 14624 2716
rect 14658 2700 14674 2734
rect 14608 2684 14674 2700
rect 14708 2726 14803 2742
rect 14708 2692 14738 2726
rect 14772 2692 14803 2726
rect 11818 2585 11849 2619
rect 11883 2585 11945 2619
rect 11979 2585 12041 2619
rect 12075 2585 12137 2619
rect 12171 2585 12233 2619
rect 12267 2585 12329 2619
rect 12363 2585 12425 2619
rect 12459 2585 12521 2619
rect 12555 2585 12617 2619
rect 12651 2585 12713 2619
rect 12747 2585 12809 2619
rect 12843 2585 12905 2619
rect 12939 2585 13001 2619
rect 13035 2585 13097 2619
rect 13131 2585 13193 2619
rect 13227 2585 13289 2619
rect 13323 2585 13385 2619
rect 13419 2585 13481 2619
rect 13515 2585 13546 2619
rect 14017 2617 14088 2648
rect 14506 2648 14522 2682
rect 14556 2648 14572 2682
rect 14506 2617 14572 2648
rect 14708 2617 14803 2692
rect 14901 2737 15156 2753
rect 14901 2703 14917 2737
rect 14951 2719 15156 2737
rect 15190 2746 15410 2762
rect 15190 2728 15360 2746
rect 14951 2703 14967 2719
rect 14901 2687 14967 2703
rect 15190 2685 15224 2728
rect 15344 2712 15360 2728
rect 15394 2712 15410 2746
rect 15344 2696 15410 2712
rect 15448 2738 15498 2754
rect 15448 2704 15464 2738
rect 15003 2651 15019 2685
rect 15053 2651 15113 2685
rect 15147 2651 15224 2685
rect 15258 2678 15308 2694
rect 15292 2644 15308 2678
rect 15258 2617 15308 2644
rect 15448 2617 15498 2704
rect 15534 2720 15600 2776
rect 15534 2686 15550 2720
rect 15584 2686 15600 2720
rect 15534 2670 15600 2686
rect 15971 2822 16005 2960
rect 16061 2938 16199 2972
rect 16370 2961 16386 2986
rect 16420 2961 16436 2995
rect 16476 3131 16526 3147
rect 16510 3097 16526 3131
rect 16570 3138 16586 3172
rect 16620 3138 16636 3172
rect 16570 3122 16636 3138
rect 16476 3088 16526 3097
rect 16674 3104 16740 3147
rect 16674 3088 16690 3104
rect 16476 3070 16690 3088
rect 16724 3070 16740 3104
rect 16476 3054 16740 3070
rect 16775 3107 16841 3245
rect 16775 3073 16791 3107
rect 16825 3073 16841 3107
rect 16775 3057 16841 3073
rect 16968 3131 17053 3147
rect 16968 3097 16984 3131
rect 17018 3097 17053 3131
rect 16476 3039 16526 3054
rect 16510 3005 16526 3039
rect 16968 3020 17053 3097
rect 16476 2989 16526 3005
rect 16267 2946 16313 2952
rect 16061 2922 16095 2938
rect 16039 2906 16095 2922
rect 16073 2872 16095 2906
rect 16267 2912 16273 2946
rect 16307 2912 16313 2946
rect 16370 2945 16436 2961
rect 16560 2986 16984 3020
rect 17018 2986 17053 3020
rect 17087 3131 17144 3147
rect 17087 3097 17103 3131
rect 17137 3097 17144 3131
rect 17087 3047 17144 3097
rect 17178 3133 17319 3245
rect 17505 3176 17571 3245
rect 17178 3099 17194 3133
rect 17228 3099 17269 3133
rect 17303 3099 17319 3133
rect 17178 3096 17319 3099
rect 17354 3146 17418 3162
rect 17354 3112 17368 3146
rect 17402 3112 17418 3146
rect 17354 3047 17418 3112
rect 17087 3013 17103 3047
rect 17137 3036 17418 3047
rect 17137 3013 17368 3036
rect 17352 3002 17368 3013
rect 17402 3002 17418 3036
rect 17352 2986 17418 3002
rect 17505 3142 17521 3176
rect 17555 3142 17571 3176
rect 17505 3093 17571 3142
rect 17505 3059 17521 3093
rect 17555 3059 17571 3093
rect 17505 3010 17571 3059
rect 16560 2955 16594 2986
rect 16267 2911 16313 2912
rect 16470 2921 16594 2955
rect 17019 2979 17053 2986
rect 16722 2946 16793 2952
rect 16470 2911 16504 2921
rect 16039 2856 16095 2872
rect 15971 2806 16027 2822
rect 15971 2772 15993 2806
rect 15971 2716 16027 2772
rect 15971 2682 15993 2716
rect 16061 2746 16095 2856
rect 16131 2890 16197 2904
rect 16131 2856 16147 2890
rect 16181 2856 16197 2890
rect 16131 2840 16197 2856
rect 16267 2895 16377 2911
rect 16267 2861 16327 2895
rect 16361 2861 16377 2895
rect 16267 2848 16377 2861
rect 16419 2895 16504 2911
rect 16419 2861 16435 2895
rect 16469 2861 16504 2895
rect 16722 2912 16753 2946
rect 16787 2912 16793 2946
rect 16722 2895 16793 2912
rect 16419 2848 16504 2861
rect 16614 2871 16680 2887
rect 16163 2814 16197 2840
rect 16614 2837 16630 2871
rect 16664 2837 16680 2871
rect 16722 2861 16738 2895
rect 16772 2861 16793 2895
rect 16939 2946 16985 2952
rect 16939 2912 16945 2946
rect 16979 2912 16985 2946
rect 17019 2945 17264 2979
rect 17505 2976 17521 3010
rect 17555 2976 17571 3010
rect 17505 2960 17571 2976
rect 17611 3176 17662 3192
rect 17645 3142 17662 3176
rect 17611 3093 17662 3142
rect 22544 3113 22573 3147
rect 22607 3113 22665 3147
rect 22699 3113 22757 3147
rect 22791 3113 22820 3147
rect 17645 3059 17662 3093
rect 17611 3010 17662 3059
rect 17645 2976 17662 3010
rect 16939 2911 16985 2912
rect 16939 2895 17082 2911
rect 16722 2848 16793 2861
rect 16830 2872 16896 2887
rect 16830 2871 16852 2872
rect 16614 2814 16680 2837
rect 16830 2837 16846 2871
rect 16886 2838 16896 2872
rect 16939 2861 17032 2895
rect 17066 2861 17082 2895
rect 16939 2851 17082 2861
rect 17116 2895 17196 2911
rect 17116 2861 17146 2895
rect 17180 2861 17196 2895
rect 17116 2860 17196 2861
rect 16880 2837 16896 2838
rect 16830 2817 16896 2837
rect 17116 2817 17150 2860
rect 17230 2826 17264 2945
rect 17314 2916 17448 2952
rect 17314 2910 17376 2916
rect 17416 2910 17448 2916
rect 17314 2876 17330 2910
rect 17364 2876 17376 2910
rect 17432 2876 17448 2910
rect 17314 2874 17376 2876
rect 17416 2874 17448 2876
rect 17314 2860 17448 2874
rect 17496 2890 17562 2906
rect 17496 2856 17512 2890
rect 17546 2856 17562 2890
rect 17496 2826 17562 2856
rect 16830 2814 17150 2817
rect 16163 2783 17150 2814
rect 17184 2792 17562 2826
rect 17611 2846 17662 2976
rect 22612 3071 22654 3113
rect 23168 3111 23197 3145
rect 23231 3111 23289 3145
rect 23323 3111 23381 3145
rect 23415 3111 23444 3145
rect 22612 3037 22620 3071
rect 22612 3003 22654 3037
rect 22612 2969 22620 3003
rect 22612 2935 22654 2969
rect 22612 2901 22620 2935
rect 22612 2885 22654 2901
rect 22688 3071 22754 3079
rect 22688 3037 22704 3071
rect 22738 3037 22754 3071
rect 22688 3003 22754 3037
rect 22688 2969 22704 3003
rect 22738 2969 22754 3003
rect 22688 2935 22754 2969
rect 22688 2901 22704 2935
rect 22738 2901 22754 2935
rect 22688 2883 22754 2901
rect 23193 3069 23239 3111
rect 23193 3035 23205 3069
rect 23193 3001 23239 3035
rect 23193 2967 23205 3001
rect 23193 2933 23239 2967
rect 23193 2899 23205 2933
rect 23193 2883 23239 2899
rect 23273 3069 23339 3077
rect 23273 3035 23289 3069
rect 23323 3035 23339 3069
rect 23273 3001 23339 3035
rect 23273 2967 23289 3001
rect 23323 2967 23339 3001
rect 23273 2933 23339 2967
rect 23273 2899 23289 2933
rect 23323 2899 23339 2933
rect 17611 2822 17616 2846
rect 17596 2808 17616 2822
rect 17658 2808 17662 2846
rect 17596 2806 17662 2808
rect 16163 2780 16896 2783
rect 17184 2749 17218 2792
rect 17596 2772 17612 2806
rect 17646 2772 17662 2806
rect 22608 2840 22674 2849
rect 22608 2802 22618 2840
rect 22608 2801 22624 2802
rect 22658 2801 22674 2840
rect 22708 2838 22754 2883
rect 23273 2881 23339 2899
rect 23373 3069 23415 3111
rect 23776 3099 23805 3133
rect 23839 3099 23897 3133
rect 23931 3099 23989 3133
rect 24023 3099 24081 3133
rect 24115 3099 24173 3133
rect 24207 3099 24236 3133
rect 23407 3035 23415 3069
rect 23373 3001 23415 3035
rect 23407 2967 23415 3001
rect 23373 2933 23415 2967
rect 23407 2899 23415 2933
rect 23373 2883 23415 2899
rect 23802 3057 23855 3099
rect 23802 3023 23821 3057
rect 23802 2989 23855 3023
rect 23802 2955 23821 2989
rect 23802 2921 23855 2955
rect 23802 2887 23821 2921
rect 22708 2804 22720 2838
rect 16061 2723 16408 2746
rect 16061 2712 16358 2723
rect 15971 2666 16027 2682
rect 16342 2689 16358 2712
rect 16392 2689 16408 2723
rect 16079 2644 16097 2678
rect 16131 2644 16150 2678
rect 16342 2667 16408 2689
rect 16450 2730 16736 2746
rect 16450 2696 16474 2730
rect 16508 2712 16686 2730
rect 16508 2696 16532 2712
rect 16450 2680 16532 2696
rect 16670 2696 16686 2712
rect 16720 2696 16736 2730
rect 16670 2680 16736 2696
rect 16770 2722 16865 2738
rect 16770 2688 16800 2722
rect 16834 2688 16865 2722
rect 13892 2583 13923 2617
rect 13957 2583 14019 2617
rect 14053 2583 14115 2617
rect 14149 2583 14211 2617
rect 14245 2583 14307 2617
rect 14341 2583 14403 2617
rect 14437 2583 14499 2617
rect 14533 2583 14595 2617
rect 14629 2583 14691 2617
rect 14725 2583 14787 2617
rect 14821 2583 14883 2617
rect 14917 2583 14979 2617
rect 15013 2583 15075 2617
rect 15109 2583 15171 2617
rect 15205 2583 15267 2617
rect 15301 2583 15363 2617
rect 15397 2583 15459 2617
rect 15493 2583 15555 2617
rect 15589 2583 15620 2617
rect 16079 2613 16150 2644
rect 16568 2644 16584 2678
rect 16618 2644 16634 2678
rect 16568 2613 16634 2644
rect 16770 2613 16865 2688
rect 16963 2733 17218 2749
rect 16963 2699 16979 2733
rect 17013 2715 17218 2733
rect 17252 2742 17472 2758
rect 17252 2724 17422 2742
rect 17013 2699 17029 2715
rect 16963 2683 17029 2699
rect 17252 2681 17286 2724
rect 17406 2708 17422 2724
rect 17456 2708 17472 2742
rect 17406 2692 17472 2708
rect 17510 2734 17560 2750
rect 17510 2700 17526 2734
rect 17065 2647 17081 2681
rect 17115 2647 17175 2681
rect 17209 2647 17286 2681
rect 17320 2674 17370 2690
rect 17354 2640 17370 2674
rect 17320 2613 17370 2640
rect 17510 2613 17560 2700
rect 17596 2716 17662 2772
rect 17596 2682 17612 2716
rect 17646 2682 17662 2716
rect 17596 2666 17662 2682
rect 22608 2751 22654 2767
rect 22708 2763 22754 2804
rect 23189 2838 23255 2849
rect 23189 2804 23196 2838
rect 23230 2833 23255 2838
rect 23189 2799 23205 2804
rect 23239 2799 23255 2833
rect 23289 2824 23339 2881
rect 23802 2871 23855 2887
rect 23889 3057 23955 3065
rect 23889 3023 23905 3057
rect 23939 3023 23955 3057
rect 23889 2989 23955 3023
rect 23889 2955 23905 2989
rect 23939 2955 23955 2989
rect 23889 2921 23955 2955
rect 23989 3057 24023 3099
rect 23989 2989 24023 3023
rect 23989 2939 24023 2955
rect 24057 3057 24123 3065
rect 24057 3023 24073 3057
rect 24107 3023 24123 3057
rect 24057 2989 24123 3023
rect 24157 3057 24199 3099
rect 24600 3085 24629 3119
rect 24663 3085 24721 3119
rect 24755 3085 24813 3119
rect 24847 3085 24905 3119
rect 24939 3085 24997 3119
rect 25031 3085 25089 3119
rect 25123 3085 25181 3119
rect 25215 3085 25244 3119
rect 24191 3023 24199 3057
rect 24157 3007 24199 3023
rect 24626 3043 24685 3085
rect 24626 3009 24635 3043
rect 24669 3009 24685 3043
rect 24057 2955 24073 2989
rect 24107 2955 24123 2989
rect 23889 2887 23905 2921
rect 23939 2905 23955 2921
rect 24057 2921 24123 2955
rect 24057 2905 24073 2921
rect 23939 2887 24073 2905
rect 24107 2909 24123 2921
rect 24626 2975 24685 3009
rect 24626 2941 24635 2975
rect 24669 2941 24685 2975
rect 24107 2887 24210 2909
rect 23889 2871 24210 2887
rect 23289 2790 23298 2824
rect 23332 2790 23339 2824
rect 22608 2717 22620 2751
rect 22608 2683 22654 2717
rect 22608 2649 22620 2683
rect 15954 2579 15985 2613
rect 16019 2579 16081 2613
rect 16115 2579 16177 2613
rect 16211 2579 16273 2613
rect 16307 2579 16369 2613
rect 16403 2579 16465 2613
rect 16499 2579 16561 2613
rect 16595 2579 16657 2613
rect 16691 2579 16753 2613
rect 16787 2579 16849 2613
rect 16883 2579 16945 2613
rect 16979 2579 17041 2613
rect 17075 2579 17137 2613
rect 17171 2579 17233 2613
rect 17267 2579 17329 2613
rect 17363 2579 17425 2613
rect 17459 2579 17521 2613
rect 17555 2579 17617 2613
rect 17651 2579 17682 2613
rect 22608 2603 22654 2649
rect 22688 2751 22754 2763
rect 22688 2717 22704 2751
rect 22738 2717 22754 2751
rect 22688 2683 22754 2717
rect 22688 2649 22704 2683
rect 22738 2649 22754 2683
rect 22688 2637 22754 2649
rect 23193 2749 23239 2765
rect 23289 2761 23339 2790
rect 23797 2822 24123 2837
rect 23797 2821 23832 2822
rect 23866 2821 24123 2822
rect 23797 2787 23813 2821
rect 23866 2788 23905 2821
rect 23847 2787 23905 2788
rect 23939 2787 23989 2821
rect 24023 2787 24073 2821
rect 24107 2787 24123 2821
rect 24157 2818 24210 2871
rect 24626 2907 24685 2941
rect 24626 2873 24635 2907
rect 24669 2873 24685 2907
rect 24626 2857 24685 2873
rect 24737 3043 24803 3051
rect 24737 3009 24753 3043
rect 24787 3009 24803 3043
rect 24737 2975 24803 3009
rect 24737 2941 24753 2975
rect 24787 2941 24803 2975
rect 24737 2907 24803 2941
rect 24837 3043 24871 3085
rect 24837 2975 24871 3009
rect 24837 2925 24871 2941
rect 24905 3043 24971 3051
rect 24905 3009 24921 3043
rect 24955 3009 24971 3043
rect 24905 2975 24971 3009
rect 24905 2941 24921 2975
rect 24955 2941 24971 2975
rect 24737 2873 24753 2907
rect 24787 2891 24803 2907
rect 24905 2907 24971 2941
rect 25005 3043 25039 3085
rect 25005 2975 25039 3009
rect 25005 2925 25039 2941
rect 25073 3043 25139 3051
rect 25073 3009 25089 3043
rect 25123 3009 25139 3043
rect 25073 2975 25139 3009
rect 25173 3043 25207 3085
rect 25173 2993 25207 3009
rect 25073 2941 25089 2975
rect 25123 2941 25139 2975
rect 24905 2891 24921 2907
rect 24787 2873 24921 2891
rect 24955 2891 24971 2907
rect 25073 2907 25139 2941
rect 25073 2891 25089 2907
rect 24955 2873 25089 2891
rect 25123 2895 25139 2907
rect 25123 2873 25227 2895
rect 24737 2857 25227 2873
rect 24157 2784 24174 2818
rect 24208 2784 24210 2818
rect 23193 2715 23205 2749
rect 23193 2677 23239 2715
rect 23193 2643 23205 2677
rect 22544 2569 22573 2603
rect 22607 2569 22665 2603
rect 22699 2569 22757 2603
rect 22791 2569 22820 2603
rect 23193 2601 23239 2643
rect 23273 2749 23339 2761
rect 23273 2715 23289 2749
rect 23323 2715 23339 2749
rect 23273 2677 23339 2715
rect 23273 2643 23289 2677
rect 23323 2643 23339 2677
rect 23273 2635 23339 2643
rect 23373 2749 23415 2765
rect 24157 2753 24210 2784
rect 24621 2814 25123 2823
rect 24621 2807 24642 2814
rect 24682 2807 25123 2814
rect 24621 2773 24637 2807
rect 24682 2776 24905 2807
rect 24671 2773 24905 2776
rect 24939 2773 24989 2807
rect 25023 2773 25073 2807
rect 25107 2773 25123 2807
rect 25157 2820 25227 2857
rect 25157 2780 25182 2820
rect 25218 2780 25227 2820
rect 23407 2715 23415 2749
rect 23373 2677 23415 2715
rect 23889 2717 24210 2753
rect 25157 2739 25227 2780
rect 23407 2643 23415 2677
rect 23373 2601 23415 2643
rect 23802 2665 23855 2681
rect 23802 2631 23821 2665
rect 23168 2567 23197 2601
rect 23231 2567 23289 2601
rect 23323 2567 23381 2601
rect 23415 2567 23444 2601
rect 23802 2589 23855 2631
rect 23889 2673 23955 2717
rect 23889 2639 23905 2673
rect 23939 2639 23955 2673
rect 23889 2623 23955 2639
rect 23989 2665 24023 2681
rect 23989 2589 24023 2631
rect 24057 2673 24123 2717
rect 24753 2703 25227 2739
rect 24057 2639 24073 2673
rect 24107 2639 24123 2673
rect 24057 2623 24123 2639
rect 24157 2666 24207 2682
rect 24191 2632 24207 2666
rect 24157 2589 24207 2632
rect 24626 2651 24679 2667
rect 24626 2617 24645 2651
rect 23776 2555 23805 2589
rect 23839 2555 23897 2589
rect 23931 2555 23989 2589
rect 24023 2555 24081 2589
rect 24115 2555 24173 2589
rect 24207 2555 24236 2589
rect 24626 2575 24679 2617
rect 24753 2659 24787 2703
rect 24753 2609 24787 2625
rect 24837 2651 24871 2667
rect 24837 2575 24871 2617
rect 24921 2659 24955 2703
rect 24921 2609 24955 2625
rect 25005 2651 25039 2667
rect 25005 2575 25039 2617
rect 25089 2659 25123 2703
rect 25089 2609 25123 2625
rect 25157 2652 25207 2668
rect 25157 2618 25173 2652
rect 25157 2575 25207 2618
rect 24600 2541 24629 2575
rect 24663 2541 24721 2575
rect 24755 2541 24813 2575
rect 24847 2541 24905 2575
rect 24939 2541 24997 2575
rect 25031 2541 25089 2575
rect 25123 2541 25181 2575
rect 25215 2541 25244 2575
<< viali >>
rect 8129 4435 8163 4469
rect 8225 4435 8259 4469
rect 8321 4435 8355 4469
rect 8220 4096 8256 4138
rect 8320 4142 8349 4146
rect 8349 4142 8354 4146
rect 8320 4112 8354 4142
rect 8129 3769 8163 3803
rect 8225 3769 8259 3803
rect 8321 3769 8355 3803
rect 1529 3269 1563 3303
rect 1625 3269 1659 3303
rect 1721 3269 1755 3303
rect 1817 3269 1851 3303
rect 1913 3269 1947 3303
rect 2009 3269 2043 3303
rect 2105 3269 2139 3303
rect 2201 3269 2235 3303
rect 2297 3269 2331 3303
rect 2393 3269 2427 3303
rect 2489 3269 2523 3303
rect 2585 3269 2619 3303
rect 2681 3269 2715 3303
rect 2777 3269 2811 3303
rect 2873 3269 2907 3303
rect 2969 3269 3003 3303
rect 3065 3269 3099 3303
rect 3161 3269 3195 3303
rect 1817 2936 1851 2970
rect 3591 3265 3625 3299
rect 3687 3265 3721 3299
rect 3783 3265 3817 3299
rect 3879 3265 3913 3299
rect 3975 3265 4009 3299
rect 4071 3265 4105 3299
rect 4167 3265 4201 3299
rect 4263 3265 4297 3299
rect 4359 3265 4393 3299
rect 4455 3265 4489 3299
rect 4551 3265 4585 3299
rect 4647 3265 4681 3299
rect 4743 3265 4777 3299
rect 4839 3265 4873 3299
rect 4935 3265 4969 3299
rect 5031 3265 5065 3299
rect 5127 3265 5161 3299
rect 5223 3265 5257 3299
rect 2297 2936 2331 2970
rect 2489 2936 2523 2970
rect 2396 2895 2430 2896
rect 2396 2862 2424 2895
rect 2424 2862 2430 2895
rect 2920 2934 2960 2940
rect 2920 2900 2942 2934
rect 2942 2900 2960 2934
rect 2920 2898 2960 2900
rect 3174 2926 3208 2960
rect 3879 2932 3913 2966
rect 5665 3263 5699 3297
rect 5761 3263 5795 3297
rect 5857 3263 5891 3297
rect 5953 3263 5987 3297
rect 6049 3263 6083 3297
rect 6145 3263 6179 3297
rect 6241 3263 6275 3297
rect 6337 3263 6371 3297
rect 6433 3263 6467 3297
rect 6529 3263 6563 3297
rect 6625 3263 6659 3297
rect 6721 3263 6755 3297
rect 6817 3263 6851 3297
rect 6913 3263 6947 3297
rect 7009 3263 7043 3297
rect 7105 3263 7139 3297
rect 7201 3263 7235 3297
rect 7297 3263 7331 3297
rect 4359 2932 4393 2966
rect 4551 2932 4585 2966
rect 4458 2891 4492 2892
rect 4458 2858 4486 2891
rect 4486 2858 4492 2891
rect 4982 2930 5022 2936
rect 4982 2896 5004 2930
rect 5004 2896 5022 2930
rect 5232 2928 5268 2962
rect 4982 2894 5022 2896
rect 1529 2603 1563 2637
rect 1625 2603 1659 2637
rect 1721 2603 1755 2637
rect 1817 2603 1851 2637
rect 1913 2603 1947 2637
rect 2009 2603 2043 2637
rect 2105 2603 2139 2637
rect 2201 2603 2235 2637
rect 2297 2603 2331 2637
rect 2393 2603 2427 2637
rect 2489 2603 2523 2637
rect 2585 2603 2619 2637
rect 2681 2603 2715 2637
rect 2777 2603 2811 2637
rect 2873 2603 2907 2637
rect 2969 2603 3003 2637
rect 3065 2603 3099 2637
rect 3161 2603 3195 2637
rect 5953 2930 5987 2964
rect 7727 3259 7761 3293
rect 7823 3259 7857 3293
rect 7919 3259 7953 3293
rect 8015 3259 8049 3293
rect 8111 3259 8145 3293
rect 8207 3259 8241 3293
rect 8303 3259 8337 3293
rect 8399 3259 8433 3293
rect 8495 3259 8529 3293
rect 8591 3259 8625 3293
rect 8687 3259 8721 3293
rect 8783 3259 8817 3293
rect 8879 3259 8913 3293
rect 8975 3259 9009 3293
rect 9071 3259 9105 3293
rect 9167 3259 9201 3293
rect 9263 3259 9297 3293
rect 9359 3259 9393 3293
rect 6433 2930 6467 2964
rect 6625 2930 6659 2964
rect 6532 2889 6566 2890
rect 6532 2856 6560 2889
rect 6560 2856 6566 2889
rect 7056 2928 7096 2934
rect 7056 2894 7078 2928
rect 7078 2894 7096 2928
rect 7056 2892 7096 2894
rect 7310 2920 7344 2954
rect 3591 2599 3625 2633
rect 3687 2599 3721 2633
rect 3783 2599 3817 2633
rect 3879 2599 3913 2633
rect 3975 2599 4009 2633
rect 4071 2599 4105 2633
rect 4167 2599 4201 2633
rect 4263 2599 4297 2633
rect 4359 2599 4393 2633
rect 4455 2599 4489 2633
rect 4551 2599 4585 2633
rect 4647 2599 4681 2633
rect 4743 2599 4777 2633
rect 4839 2599 4873 2633
rect 4935 2599 4969 2633
rect 5031 2599 5065 2633
rect 5127 2599 5161 2633
rect 5223 2599 5257 2633
rect 8015 2926 8049 2960
rect 9787 3255 9821 3289
rect 9883 3255 9917 3289
rect 9979 3255 10013 3289
rect 10075 3255 10109 3289
rect 10171 3255 10205 3289
rect 10267 3255 10301 3289
rect 10363 3255 10397 3289
rect 10459 3255 10493 3289
rect 10555 3255 10589 3289
rect 10651 3255 10685 3289
rect 10747 3255 10781 3289
rect 10843 3255 10877 3289
rect 10939 3255 10973 3289
rect 11035 3255 11069 3289
rect 11131 3255 11165 3289
rect 11227 3255 11261 3289
rect 11323 3255 11357 3289
rect 11419 3255 11453 3289
rect 8495 2926 8529 2960
rect 8687 2926 8721 2960
rect 8594 2885 8628 2886
rect 8594 2852 8622 2885
rect 8622 2852 8628 2885
rect 9118 2924 9158 2930
rect 9118 2890 9140 2924
rect 9140 2890 9158 2924
rect 9118 2888 9158 2890
rect 9366 2910 9402 2944
rect 5665 2597 5699 2631
rect 5761 2597 5795 2631
rect 5857 2597 5891 2631
rect 5953 2597 5987 2631
rect 6049 2597 6083 2631
rect 6145 2597 6179 2631
rect 6241 2597 6275 2631
rect 6337 2597 6371 2631
rect 6433 2597 6467 2631
rect 6529 2597 6563 2631
rect 6625 2597 6659 2631
rect 6721 2597 6755 2631
rect 6817 2597 6851 2631
rect 6913 2597 6947 2631
rect 7009 2597 7043 2631
rect 7105 2597 7139 2631
rect 7201 2597 7235 2631
rect 7297 2597 7331 2631
rect 10075 2922 10109 2956
rect 11849 3251 11883 3285
rect 11945 3251 11979 3285
rect 12041 3251 12075 3285
rect 12137 3251 12171 3285
rect 12233 3251 12267 3285
rect 12329 3251 12363 3285
rect 12425 3251 12459 3285
rect 12521 3251 12555 3285
rect 12617 3251 12651 3285
rect 12713 3251 12747 3285
rect 12809 3251 12843 3285
rect 12905 3251 12939 3285
rect 13001 3251 13035 3285
rect 13097 3251 13131 3285
rect 13193 3251 13227 3285
rect 13289 3251 13323 3285
rect 13385 3251 13419 3285
rect 13481 3251 13515 3285
rect 10555 2922 10589 2956
rect 10747 2922 10781 2956
rect 10654 2881 10688 2882
rect 10654 2848 10682 2881
rect 10682 2848 10688 2881
rect 11178 2920 11218 2926
rect 11178 2886 11200 2920
rect 11200 2886 11218 2920
rect 11178 2884 11218 2886
rect 11432 2912 11466 2946
rect 7727 2593 7761 2627
rect 7823 2593 7857 2627
rect 7919 2593 7953 2627
rect 8015 2593 8049 2627
rect 8111 2593 8145 2627
rect 8207 2593 8241 2627
rect 8303 2593 8337 2627
rect 8399 2593 8433 2627
rect 8495 2593 8529 2627
rect 8591 2593 8625 2627
rect 8687 2593 8721 2627
rect 8783 2593 8817 2627
rect 8879 2593 8913 2627
rect 8975 2593 9009 2627
rect 9071 2593 9105 2627
rect 9167 2593 9201 2627
rect 9263 2593 9297 2627
rect 9359 2593 9393 2627
rect 12137 2918 12171 2952
rect 13923 3249 13957 3283
rect 14019 3249 14053 3283
rect 14115 3249 14149 3283
rect 14211 3249 14245 3283
rect 14307 3249 14341 3283
rect 14403 3249 14437 3283
rect 14499 3249 14533 3283
rect 14595 3249 14629 3283
rect 14691 3249 14725 3283
rect 14787 3249 14821 3283
rect 14883 3249 14917 3283
rect 14979 3249 15013 3283
rect 15075 3249 15109 3283
rect 15171 3249 15205 3283
rect 15267 3249 15301 3283
rect 15363 3249 15397 3283
rect 15459 3249 15493 3283
rect 15555 3249 15589 3283
rect 12617 2918 12651 2952
rect 12809 2918 12843 2952
rect 12716 2877 12750 2878
rect 12716 2844 12744 2877
rect 12744 2844 12750 2877
rect 13240 2916 13280 2922
rect 13240 2882 13262 2916
rect 13262 2882 13280 2916
rect 13490 2914 13526 2948
rect 13240 2880 13280 2882
rect 9787 2589 9821 2623
rect 9883 2589 9917 2623
rect 9979 2589 10013 2623
rect 10075 2589 10109 2623
rect 10171 2589 10205 2623
rect 10267 2589 10301 2623
rect 10363 2589 10397 2623
rect 10459 2589 10493 2623
rect 10555 2589 10589 2623
rect 10651 2589 10685 2623
rect 10747 2589 10781 2623
rect 10843 2589 10877 2623
rect 10939 2589 10973 2623
rect 11035 2589 11069 2623
rect 11131 2589 11165 2623
rect 11227 2589 11261 2623
rect 11323 2589 11357 2623
rect 11419 2589 11453 2623
rect 14211 2916 14245 2950
rect 15985 3245 16019 3279
rect 16081 3245 16115 3279
rect 16177 3245 16211 3279
rect 16273 3245 16307 3279
rect 16369 3245 16403 3279
rect 16465 3245 16499 3279
rect 16561 3245 16595 3279
rect 16657 3245 16691 3279
rect 16753 3245 16787 3279
rect 16849 3245 16883 3279
rect 16945 3245 16979 3279
rect 17041 3245 17075 3279
rect 17137 3245 17171 3279
rect 17233 3245 17267 3279
rect 17329 3245 17363 3279
rect 17425 3245 17459 3279
rect 17521 3245 17555 3279
rect 17617 3245 17651 3279
rect 14691 2916 14725 2950
rect 14883 2916 14917 2950
rect 14790 2875 14824 2876
rect 14790 2842 14818 2875
rect 14818 2842 14824 2875
rect 15314 2914 15354 2920
rect 15314 2880 15336 2914
rect 15336 2880 15354 2914
rect 15314 2878 15354 2880
rect 15568 2906 15602 2940
rect 11849 2585 11883 2619
rect 11945 2585 11979 2619
rect 12041 2585 12075 2619
rect 12137 2585 12171 2619
rect 12233 2585 12267 2619
rect 12329 2585 12363 2619
rect 12425 2585 12459 2619
rect 12521 2585 12555 2619
rect 12617 2585 12651 2619
rect 12713 2585 12747 2619
rect 12809 2585 12843 2619
rect 12905 2585 12939 2619
rect 13001 2585 13035 2619
rect 13097 2585 13131 2619
rect 13193 2585 13227 2619
rect 13289 2585 13323 2619
rect 13385 2585 13419 2619
rect 13481 2585 13515 2619
rect 16273 2912 16307 2946
rect 16753 2912 16787 2946
rect 16945 2912 16979 2946
rect 22573 3113 22607 3147
rect 22665 3113 22699 3147
rect 22757 3113 22791 3147
rect 16852 2871 16886 2872
rect 16852 2838 16880 2871
rect 16880 2838 16886 2871
rect 17376 2910 17416 2916
rect 17376 2876 17398 2910
rect 17398 2876 17416 2910
rect 17376 2874 17416 2876
rect 23197 3111 23231 3145
rect 23289 3111 23323 3145
rect 23381 3111 23415 3145
rect 17616 2808 17658 2846
rect 22618 2835 22658 2840
rect 22618 2802 22624 2835
rect 22624 2802 22658 2835
rect 23805 3099 23839 3133
rect 23897 3099 23931 3133
rect 23989 3099 24023 3133
rect 24081 3099 24115 3133
rect 24173 3099 24207 3133
rect 22720 2804 22754 2838
rect 13923 2583 13957 2617
rect 14019 2583 14053 2617
rect 14115 2583 14149 2617
rect 14211 2583 14245 2617
rect 14307 2583 14341 2617
rect 14403 2583 14437 2617
rect 14499 2583 14533 2617
rect 14595 2583 14629 2617
rect 14691 2583 14725 2617
rect 14787 2583 14821 2617
rect 14883 2583 14917 2617
rect 14979 2583 15013 2617
rect 15075 2583 15109 2617
rect 15171 2583 15205 2617
rect 15267 2583 15301 2617
rect 15363 2583 15397 2617
rect 15459 2583 15493 2617
rect 15555 2583 15589 2617
rect 23196 2833 23230 2838
rect 23196 2804 23205 2833
rect 23205 2804 23230 2833
rect 24629 3085 24663 3119
rect 24721 3085 24755 3119
rect 24813 3085 24847 3119
rect 24905 3085 24939 3119
rect 24997 3085 25031 3119
rect 25089 3085 25123 3119
rect 25181 3085 25215 3119
rect 23298 2790 23332 2824
rect 15985 2579 16019 2613
rect 16081 2579 16115 2613
rect 16177 2579 16211 2613
rect 16273 2579 16307 2613
rect 16369 2579 16403 2613
rect 16465 2579 16499 2613
rect 16561 2579 16595 2613
rect 16657 2579 16691 2613
rect 16753 2579 16787 2613
rect 16849 2579 16883 2613
rect 16945 2579 16979 2613
rect 17041 2579 17075 2613
rect 17137 2579 17171 2613
rect 17233 2579 17267 2613
rect 17329 2579 17363 2613
rect 17425 2579 17459 2613
rect 17521 2579 17555 2613
rect 17617 2579 17651 2613
rect 23832 2821 23866 2822
rect 23832 2788 23847 2821
rect 23847 2788 23866 2821
rect 24174 2784 24208 2818
rect 22573 2569 22607 2603
rect 22665 2569 22699 2603
rect 22757 2569 22791 2603
rect 24642 2807 24682 2814
rect 24642 2776 24671 2807
rect 24671 2776 24682 2807
rect 25182 2780 25218 2820
rect 23197 2567 23231 2601
rect 23289 2567 23323 2601
rect 23381 2567 23415 2601
rect 23805 2555 23839 2589
rect 23897 2555 23931 2589
rect 23989 2555 24023 2589
rect 24081 2555 24115 2589
rect 24173 2555 24207 2589
rect 24629 2541 24663 2575
rect 24721 2541 24755 2575
rect 24813 2541 24847 2575
rect 24905 2541 24939 2575
rect 24997 2541 25031 2575
rect 25089 2541 25123 2575
rect 25181 2541 25215 2575
<< metal1 >>
rect 890 4486 972 4516
rect 890 4420 904 4486
rect 958 4473 972 4486
rect 8098 4473 8386 4501
rect 958 4469 8386 4473
rect 958 4441 8129 4469
rect 958 4420 972 4441
rect 890 4386 972 4420
rect 8098 4435 8129 4441
rect 8163 4435 8225 4469
rect 8259 4435 8321 4469
rect 8355 4435 8386 4469
rect 8098 4403 8386 4435
rect 8182 4142 8266 4174
rect 17763 4172 17869 4181
rect 8182 4090 8192 4142
rect 8244 4138 8266 4142
rect 8256 4096 8266 4138
rect 8244 4090 8266 4096
rect 8182 4060 8266 4090
rect 8307 4146 17869 4172
rect 8307 4112 8320 4146
rect 8354 4112 17869 4146
rect 8307 4086 17869 4112
rect 8220 4044 8265 4060
rect 294 3830 484 3880
rect 294 3740 344 3830
rect 438 3807 484 3830
rect 8098 3807 8386 3835
rect 438 3803 8386 3807
rect 438 3775 8129 3803
rect 438 3740 484 3775
rect 294 3684 484 3740
rect 8098 3769 8129 3775
rect 8163 3769 8225 3803
rect 8259 3769 8321 3803
rect 8355 3769 8386 3803
rect 8098 3737 8386 3769
rect 354 3322 466 3390
rect 1498 3322 3226 3335
rect 354 3320 3226 3322
rect 354 3228 366 3320
rect 442 3308 3226 3320
rect 3560 3308 5288 3331
rect 442 3303 5288 3308
rect 442 3269 1529 3303
rect 1563 3269 1625 3303
rect 1659 3269 1721 3303
rect 1755 3269 1817 3303
rect 1851 3269 1913 3303
rect 1947 3269 2009 3303
rect 2043 3269 2105 3303
rect 2139 3269 2201 3303
rect 2235 3269 2297 3303
rect 2331 3269 2393 3303
rect 2427 3269 2489 3303
rect 2523 3269 2585 3303
rect 2619 3269 2681 3303
rect 2715 3269 2777 3303
rect 2811 3269 2873 3303
rect 2907 3269 2969 3303
rect 3003 3269 3065 3303
rect 3099 3269 3161 3303
rect 3195 3299 5288 3303
rect 3195 3269 3591 3299
rect 442 3265 3591 3269
rect 3625 3265 3687 3299
rect 3721 3265 3783 3299
rect 3817 3265 3879 3299
rect 3913 3265 3975 3299
rect 4009 3265 4071 3299
rect 4105 3265 4167 3299
rect 4201 3265 4263 3299
rect 4297 3265 4359 3299
rect 4393 3265 4455 3299
rect 4489 3265 4551 3299
rect 4585 3265 4647 3299
rect 4681 3265 4743 3299
rect 4777 3265 4839 3299
rect 4873 3265 4935 3299
rect 4969 3265 5031 3299
rect 5065 3265 5127 3299
rect 5161 3265 5223 3299
rect 5257 3298 5288 3299
rect 5634 3298 7362 3329
rect 7696 3300 9424 3325
rect 9756 3300 11484 3321
rect 7696 3298 11484 3300
rect 5257 3297 11484 3298
rect 5257 3265 5665 3297
rect 442 3263 5665 3265
rect 5699 3263 5761 3297
rect 5795 3263 5857 3297
rect 5891 3263 5953 3297
rect 5987 3263 6049 3297
rect 6083 3263 6145 3297
rect 6179 3263 6241 3297
rect 6275 3263 6337 3297
rect 6371 3263 6433 3297
rect 6467 3263 6529 3297
rect 6563 3263 6625 3297
rect 6659 3263 6721 3297
rect 6755 3263 6817 3297
rect 6851 3263 6913 3297
rect 6947 3263 7009 3297
rect 7043 3263 7105 3297
rect 7139 3263 7201 3297
rect 7235 3263 7297 3297
rect 7331 3293 11484 3297
rect 7331 3263 7727 3293
rect 442 3260 7727 3263
rect 442 3237 3226 3260
rect 3560 3259 7727 3260
rect 7761 3259 7823 3293
rect 7857 3259 7919 3293
rect 7953 3259 8015 3293
rect 8049 3259 8111 3293
rect 8145 3259 8207 3293
rect 8241 3259 8303 3293
rect 8337 3259 8399 3293
rect 8433 3259 8495 3293
rect 8529 3259 8591 3293
rect 8625 3259 8687 3293
rect 8721 3259 8783 3293
rect 8817 3259 8879 3293
rect 8913 3259 8975 3293
rect 9009 3259 9071 3293
rect 9105 3259 9167 3293
rect 9201 3259 9263 3293
rect 9297 3259 9359 3293
rect 9393 3289 11484 3293
rect 9393 3259 9787 3289
rect 3560 3255 9787 3259
rect 9821 3255 9883 3289
rect 9917 3255 9979 3289
rect 10013 3255 10075 3289
rect 10109 3255 10171 3289
rect 10205 3255 10267 3289
rect 10301 3255 10363 3289
rect 10397 3255 10459 3289
rect 10493 3255 10555 3289
rect 10589 3255 10651 3289
rect 10685 3255 10747 3289
rect 10781 3255 10843 3289
rect 10877 3255 10939 3289
rect 10973 3255 11035 3289
rect 11069 3255 11131 3289
rect 11165 3255 11227 3289
rect 11261 3255 11323 3289
rect 11357 3255 11419 3289
rect 11453 3286 11484 3289
rect 11818 3290 13546 3317
rect 13892 3290 15620 3315
rect 15954 3290 17682 3311
rect 11818 3286 17682 3290
rect 11453 3285 17682 3286
rect 11453 3255 11849 3285
rect 3560 3252 11849 3255
rect 3560 3250 9424 3252
rect 442 3236 1604 3237
rect 442 3228 466 3236
rect 354 3166 466 3228
rect 2096 2988 2192 3010
rect 1805 2970 1863 2976
rect 1805 2936 1817 2970
rect 1851 2967 1863 2970
rect 2096 2967 2132 2988
rect 1851 2939 2132 2967
rect 1851 2936 1863 2939
rect 1805 2930 1863 2936
rect 2096 2936 2132 2939
rect 2184 2967 2192 2988
rect 2285 2970 2343 2976
rect 2285 2967 2297 2970
rect 2184 2939 2297 2967
rect 2184 2936 2192 2939
rect 2096 2910 2192 2936
rect 2285 2936 2297 2939
rect 2331 2967 2343 2970
rect 2477 2970 2535 2976
rect 2918 2974 2972 3237
rect 3560 3233 5288 3250
rect 2477 2967 2489 2970
rect 2331 2939 2489 2967
rect 2331 2936 2343 2939
rect 2285 2930 2343 2936
rect 2477 2936 2489 2939
rect 2523 2936 2535 2970
rect 2477 2930 2535 2936
rect 2858 2940 2990 2974
rect 2376 2896 2446 2910
rect 2376 2862 2396 2896
rect 2430 2862 2446 2896
rect 2858 2898 2920 2940
rect 2960 2898 2990 2940
rect 3166 2972 3920 2978
rect 3166 2966 3925 2972
rect 3166 2960 3879 2966
rect 3166 2926 3174 2960
rect 3208 2932 3879 2960
rect 3913 2963 3925 2966
rect 4347 2966 4405 2972
rect 4347 2963 4359 2966
rect 3913 2935 4359 2963
rect 3913 2932 3925 2935
rect 3208 2926 3925 2932
rect 4347 2932 4359 2935
rect 4393 2963 4405 2966
rect 4539 2966 4597 2972
rect 4980 2970 5034 3233
rect 5634 3231 7362 3250
rect 5218 2972 5274 3004
rect 5218 2970 5978 2972
rect 4539 2963 4551 2966
rect 4393 2935 4551 2963
rect 4393 2932 4405 2935
rect 4347 2926 4405 2932
rect 4539 2932 4551 2935
rect 4585 2932 4597 2966
rect 4539 2926 4597 2932
rect 4920 2936 5052 2970
rect 3166 2912 3920 2926
rect 2858 2888 2990 2898
rect 4438 2892 4508 2906
rect 2376 2830 2446 2862
rect 4438 2858 4458 2892
rect 4492 2858 4508 2892
rect 4920 2894 4982 2936
rect 5022 2894 5052 2936
rect 5218 2964 5999 2970
rect 5218 2962 5953 2964
rect 5218 2928 5232 2962
rect 5268 2930 5953 2962
rect 5987 2961 5999 2964
rect 6421 2964 6479 2970
rect 6421 2961 6433 2964
rect 5987 2933 6433 2961
rect 5987 2930 5999 2933
rect 5268 2928 5999 2930
rect 5218 2924 5999 2928
rect 6421 2930 6433 2933
rect 6467 2961 6479 2964
rect 6613 2964 6671 2970
rect 7054 2968 7108 3231
rect 7696 3227 9424 3250
rect 9756 3251 11849 3252
rect 11883 3251 11945 3285
rect 11979 3251 12041 3285
rect 12075 3251 12137 3285
rect 12171 3251 12233 3285
rect 12267 3251 12329 3285
rect 12363 3251 12425 3285
rect 12459 3251 12521 3285
rect 12555 3251 12617 3285
rect 12651 3251 12713 3285
rect 12747 3251 12809 3285
rect 12843 3251 12905 3285
rect 12939 3251 13001 3285
rect 13035 3251 13097 3285
rect 13131 3251 13193 3285
rect 13227 3251 13289 3285
rect 13323 3251 13385 3285
rect 13419 3251 13481 3285
rect 13515 3283 17682 3285
rect 13515 3251 13923 3283
rect 9756 3249 13923 3251
rect 13957 3249 14019 3283
rect 14053 3249 14115 3283
rect 14149 3249 14211 3283
rect 14245 3249 14307 3283
rect 14341 3249 14403 3283
rect 14437 3249 14499 3283
rect 14533 3249 14595 3283
rect 14629 3249 14691 3283
rect 14725 3249 14787 3283
rect 14821 3249 14883 3283
rect 14917 3249 14979 3283
rect 15013 3249 15075 3283
rect 15109 3249 15171 3283
rect 15205 3249 15267 3283
rect 15301 3249 15363 3283
rect 15397 3249 15459 3283
rect 15493 3249 15555 3283
rect 15589 3279 17682 3283
rect 15589 3249 15985 3279
rect 9756 3245 15985 3249
rect 16019 3245 16081 3279
rect 16115 3245 16177 3279
rect 16211 3245 16273 3279
rect 16307 3245 16369 3279
rect 16403 3245 16465 3279
rect 16499 3245 16561 3279
rect 16595 3245 16657 3279
rect 16691 3245 16753 3279
rect 16787 3245 16849 3279
rect 16883 3245 16945 3279
rect 16979 3245 17041 3279
rect 17075 3245 17137 3279
rect 17171 3245 17233 3279
rect 17267 3245 17329 3279
rect 17363 3245 17425 3279
rect 17459 3245 17521 3279
rect 17555 3245 17617 3279
rect 17651 3245 17682 3279
rect 9756 3242 17682 3245
rect 9756 3238 13546 3242
rect 6613 2961 6625 2964
rect 6467 2933 6625 2961
rect 6467 2930 6479 2933
rect 6421 2924 6479 2930
rect 6613 2930 6625 2933
rect 6659 2930 6671 2964
rect 6613 2924 6671 2930
rect 6994 2934 7126 2968
rect 5218 2914 5978 2924
rect 5218 2910 5274 2914
rect 4920 2884 5052 2894
rect 6512 2890 6582 2904
rect 966 2664 1096 2704
rect 2392 2669 2424 2830
rect 4438 2826 4508 2858
rect 6512 2856 6532 2890
rect 6566 2856 6582 2890
rect 6994 2892 7056 2934
rect 7096 2892 7126 2934
rect 7302 2966 8056 2972
rect 7302 2960 8061 2966
rect 7302 2954 8015 2960
rect 7302 2920 7310 2954
rect 7344 2926 8015 2954
rect 8049 2957 8061 2960
rect 8483 2960 8541 2966
rect 8483 2957 8495 2960
rect 8049 2929 8495 2957
rect 8049 2926 8061 2929
rect 7344 2920 8061 2926
rect 8483 2926 8495 2929
rect 8529 2957 8541 2960
rect 8675 2960 8733 2966
rect 9116 2964 9170 3227
rect 9756 3223 11484 3238
rect 8675 2957 8687 2960
rect 8529 2929 8687 2957
rect 8529 2926 8541 2929
rect 8483 2920 8541 2926
rect 8675 2926 8687 2929
rect 8721 2926 8733 2960
rect 8675 2920 8733 2926
rect 9056 2930 9188 2964
rect 9362 2962 10114 2966
rect 7302 2906 8056 2920
rect 6994 2882 7126 2892
rect 8574 2886 8644 2900
rect 1498 2664 3226 2669
rect 4454 2665 4486 2826
rect 6512 2824 6582 2856
rect 8574 2852 8594 2886
rect 8628 2852 8644 2886
rect 9056 2888 9118 2930
rect 9158 2888 9188 2930
rect 9354 2956 10121 2962
rect 9354 2944 10075 2956
rect 9354 2910 9366 2944
rect 9402 2922 10075 2944
rect 10109 2953 10121 2956
rect 10543 2956 10601 2962
rect 10543 2953 10555 2956
rect 10109 2925 10555 2953
rect 10109 2922 10121 2925
rect 9402 2916 10121 2922
rect 10543 2922 10555 2925
rect 10589 2953 10601 2956
rect 10735 2956 10793 2962
rect 11176 2960 11230 3223
rect 11818 3219 13546 3238
rect 10735 2953 10747 2956
rect 10589 2925 10747 2953
rect 10589 2922 10601 2925
rect 10543 2916 10601 2922
rect 10735 2922 10747 2925
rect 10781 2922 10793 2956
rect 10735 2916 10793 2922
rect 11116 2926 11248 2960
rect 9402 2910 10114 2916
rect 9354 2900 10114 2910
rect 9362 2898 10114 2900
rect 9056 2878 9188 2888
rect 10634 2882 10704 2896
rect 966 2660 3226 2664
rect 966 2582 1000 2660
rect 1066 2638 3226 2660
rect 3560 2642 5288 2665
rect 6528 2663 6560 2824
rect 8574 2820 8644 2852
rect 10634 2848 10654 2882
rect 10688 2848 10704 2882
rect 11116 2884 11178 2926
rect 11218 2884 11248 2926
rect 11424 2958 12178 2964
rect 11424 2952 12183 2958
rect 11424 2946 12137 2952
rect 11424 2912 11432 2946
rect 11466 2918 12137 2946
rect 12171 2949 12183 2952
rect 12605 2952 12663 2958
rect 12605 2949 12617 2952
rect 12171 2921 12617 2949
rect 12171 2918 12183 2921
rect 11466 2912 12183 2918
rect 12605 2918 12617 2921
rect 12651 2949 12663 2952
rect 12797 2952 12855 2958
rect 13238 2956 13292 3219
rect 13892 3217 15620 3242
rect 13476 2958 13532 2990
rect 13476 2956 14236 2958
rect 12797 2949 12809 2952
rect 12651 2921 12809 2949
rect 12651 2918 12663 2921
rect 12605 2912 12663 2918
rect 12797 2918 12809 2921
rect 12843 2918 12855 2952
rect 12797 2912 12855 2918
rect 13178 2922 13310 2956
rect 11424 2898 12178 2912
rect 11116 2874 11248 2884
rect 12696 2878 12766 2892
rect 5634 2642 7362 2663
rect 8590 2659 8622 2820
rect 10634 2816 10704 2848
rect 12696 2844 12716 2878
rect 12750 2844 12766 2878
rect 13178 2880 13240 2922
rect 13280 2880 13310 2922
rect 13476 2950 14257 2956
rect 13476 2948 14211 2950
rect 13476 2914 13490 2948
rect 13526 2916 14211 2948
rect 14245 2947 14257 2950
rect 14679 2950 14737 2956
rect 14679 2947 14691 2950
rect 14245 2919 14691 2947
rect 14245 2916 14257 2919
rect 13526 2914 14257 2916
rect 13476 2910 14257 2914
rect 14679 2916 14691 2919
rect 14725 2947 14737 2950
rect 14871 2950 14929 2956
rect 15312 2954 15366 3217
rect 15954 3213 17682 3242
rect 14871 2947 14883 2950
rect 14725 2919 14883 2947
rect 14725 2916 14737 2919
rect 14679 2910 14737 2916
rect 14871 2916 14883 2919
rect 14917 2916 14929 2950
rect 14871 2910 14929 2916
rect 15252 2920 15384 2954
rect 13476 2900 14236 2910
rect 13476 2896 13532 2900
rect 13178 2870 13310 2880
rect 14770 2876 14840 2890
rect 3560 2638 7362 2642
rect 1066 2637 7362 2638
rect 1066 2603 1529 2637
rect 1563 2603 1625 2637
rect 1659 2603 1721 2637
rect 1755 2603 1817 2637
rect 1851 2603 1913 2637
rect 1947 2603 2009 2637
rect 2043 2603 2105 2637
rect 2139 2603 2201 2637
rect 2235 2603 2297 2637
rect 2331 2603 2393 2637
rect 2427 2603 2489 2637
rect 2523 2603 2585 2637
rect 2619 2603 2681 2637
rect 2715 2603 2777 2637
rect 2811 2603 2873 2637
rect 2907 2603 2969 2637
rect 3003 2603 3065 2637
rect 3099 2603 3161 2637
rect 3195 2633 7362 2637
rect 3195 2603 3591 2633
rect 1066 2599 3591 2603
rect 3625 2599 3687 2633
rect 3721 2599 3783 2633
rect 3817 2599 3879 2633
rect 3913 2599 3975 2633
rect 4009 2599 4071 2633
rect 4105 2599 4167 2633
rect 4201 2599 4263 2633
rect 4297 2599 4359 2633
rect 4393 2599 4455 2633
rect 4489 2599 4551 2633
rect 4585 2599 4647 2633
rect 4681 2599 4743 2633
rect 4777 2599 4839 2633
rect 4873 2599 4935 2633
rect 4969 2599 5031 2633
rect 5065 2599 5127 2633
rect 5161 2599 5223 2633
rect 5257 2631 7362 2633
rect 5257 2599 5665 2631
rect 1066 2597 5665 2599
rect 5699 2597 5761 2631
rect 5795 2597 5857 2631
rect 5891 2597 5953 2631
rect 5987 2597 6049 2631
rect 6083 2597 6145 2631
rect 6179 2597 6241 2631
rect 6275 2597 6337 2631
rect 6371 2597 6433 2631
rect 6467 2597 6529 2631
rect 6563 2597 6625 2631
rect 6659 2597 6721 2631
rect 6755 2597 6817 2631
rect 6851 2597 6913 2631
rect 6947 2597 7009 2631
rect 7043 2597 7105 2631
rect 7139 2597 7201 2631
rect 7235 2597 7297 2631
rect 7331 2626 7362 2631
rect 7696 2627 9424 2659
rect 10650 2655 10682 2816
rect 12696 2812 12766 2844
rect 14770 2842 14790 2876
rect 14824 2842 14840 2876
rect 15252 2878 15314 2920
rect 15354 2878 15384 2920
rect 15560 2952 16314 2958
rect 15560 2946 16319 2952
rect 15560 2940 16273 2946
rect 15560 2906 15568 2940
rect 15602 2912 16273 2940
rect 16307 2943 16319 2946
rect 16741 2946 16799 2952
rect 16741 2943 16753 2946
rect 16307 2915 16753 2943
rect 16307 2912 16319 2915
rect 15602 2906 16319 2912
rect 16741 2912 16753 2915
rect 16787 2943 16799 2946
rect 16933 2946 16991 2952
rect 17374 2950 17428 3213
rect 16933 2943 16945 2946
rect 16787 2915 16945 2943
rect 16787 2912 16799 2915
rect 16741 2906 16799 2912
rect 16933 2912 16945 2915
rect 16979 2912 16991 2946
rect 16933 2906 16991 2912
rect 17314 2916 17446 2950
rect 15560 2892 16314 2906
rect 15252 2868 15384 2878
rect 16832 2872 16902 2886
rect 7696 2626 7727 2627
rect 7331 2597 7727 2626
rect 1066 2594 7727 2597
rect 1066 2590 5288 2594
rect 1066 2582 3226 2590
rect 966 2522 1096 2582
rect 1498 2571 3226 2582
rect 3560 2567 5288 2590
rect 5634 2593 7727 2594
rect 7761 2593 7823 2627
rect 7857 2593 7919 2627
rect 7953 2593 8015 2627
rect 8049 2593 8111 2627
rect 8145 2593 8207 2627
rect 8241 2593 8303 2627
rect 8337 2593 8399 2627
rect 8433 2593 8495 2627
rect 8529 2593 8591 2627
rect 8625 2593 8687 2627
rect 8721 2593 8783 2627
rect 8817 2593 8879 2627
rect 8913 2593 8975 2627
rect 9009 2593 9071 2627
rect 9105 2593 9167 2627
rect 9201 2593 9263 2627
rect 9297 2593 9359 2627
rect 9393 2626 9424 2627
rect 9756 2626 11484 2655
rect 12712 2651 12744 2812
rect 14770 2810 14840 2842
rect 16832 2838 16852 2872
rect 16886 2838 16902 2872
rect 17314 2874 17376 2916
rect 17416 2874 17446 2916
rect 17763 2876 17869 4086
rect 22544 3158 22820 3178
rect 22544 3147 22654 3158
rect 22706 3147 22820 3158
rect 22544 3113 22573 3147
rect 22607 3113 22654 3147
rect 22706 3113 22757 3147
rect 22791 3113 22820 3147
rect 22544 3106 22654 3113
rect 22706 3106 22820 3113
rect 22544 3082 22820 3106
rect 23168 3152 23444 3176
rect 23168 3145 23268 3152
rect 23326 3145 23444 3152
rect 23168 3111 23197 3145
rect 23231 3111 23268 3145
rect 23326 3111 23381 3145
rect 23415 3111 23444 3145
rect 23168 3096 23268 3111
rect 23326 3096 23444 3111
rect 23168 3080 23444 3096
rect 23776 3152 24236 3164
rect 23776 3133 23982 3152
rect 24040 3133 24236 3152
rect 23776 3099 23805 3133
rect 23839 3099 23897 3133
rect 23931 3099 23982 3133
rect 24040 3099 24081 3133
rect 24115 3099 24173 3133
rect 24207 3099 24236 3133
rect 23776 3096 23982 3099
rect 24040 3096 24236 3099
rect 23776 3068 24236 3096
rect 24600 3138 25244 3150
rect 24600 3119 24914 3138
rect 24972 3119 25244 3138
rect 24600 3085 24629 3119
rect 24663 3085 24721 3119
rect 24755 3085 24813 3119
rect 24847 3085 24905 3119
rect 24972 3085 24997 3119
rect 25031 3085 25089 3119
rect 25123 3085 25181 3119
rect 25215 3085 25244 3119
rect 24600 3082 24914 3085
rect 24972 3082 25244 3085
rect 24600 3054 25244 3082
rect 17314 2864 17446 2874
rect 9393 2623 11484 2626
rect 9393 2593 9787 2623
rect 5634 2589 9787 2593
rect 9821 2589 9883 2623
rect 9917 2589 9979 2623
rect 10013 2589 10075 2623
rect 10109 2589 10171 2623
rect 10205 2589 10267 2623
rect 10301 2589 10363 2623
rect 10397 2589 10459 2623
rect 10493 2589 10555 2623
rect 10589 2589 10651 2623
rect 10685 2589 10747 2623
rect 10781 2589 10843 2623
rect 10877 2589 10939 2623
rect 10973 2589 11035 2623
rect 11069 2589 11131 2623
rect 11165 2589 11227 2623
rect 11261 2589 11323 2623
rect 11357 2589 11419 2623
rect 11453 2622 11484 2623
rect 11818 2622 13546 2651
rect 14786 2649 14818 2810
rect 16832 2806 16902 2838
rect 17610 2846 22675 2876
rect 17610 2808 17616 2846
rect 17658 2840 22675 2846
rect 17658 2808 22618 2840
rect 13892 2626 15620 2649
rect 16848 2645 16880 2806
rect 17610 2802 22618 2808
rect 22658 2802 22675 2840
rect 17610 2758 22675 2802
rect 22712 2838 23258 2858
rect 22712 2804 22720 2838
rect 22754 2804 23196 2838
rect 23230 2804 23258 2838
rect 22712 2786 23258 2804
rect 23288 2826 23344 2838
rect 23796 2826 23904 2854
rect 23288 2824 23904 2826
rect 23288 2790 23298 2824
rect 23332 2822 23904 2824
rect 23332 2790 23832 2822
rect 23288 2774 23344 2790
rect 23796 2788 23832 2790
rect 23866 2788 23904 2822
rect 24158 2818 24216 2830
rect 24618 2818 24694 2846
rect 25171 2820 30510 2876
rect 23796 2776 23904 2788
rect 24156 2784 24174 2818
rect 24208 2814 24718 2818
rect 24208 2784 24642 2814
rect 24156 2776 24642 2784
rect 24682 2776 24718 2814
rect 25171 2780 25182 2820
rect 25218 2780 30510 2820
rect 24158 2770 24216 2776
rect 24618 2756 24694 2776
rect 25171 2758 30510 2780
rect 15954 2626 17682 2645
rect 13892 2622 17682 2626
rect 11453 2619 17682 2622
rect 11453 2589 11849 2619
rect 5634 2585 11849 2589
rect 11883 2585 11945 2619
rect 11979 2585 12041 2619
rect 12075 2585 12137 2619
rect 12171 2585 12233 2619
rect 12267 2585 12329 2619
rect 12363 2585 12425 2619
rect 12459 2585 12521 2619
rect 12555 2585 12617 2619
rect 12651 2585 12713 2619
rect 12747 2585 12809 2619
rect 12843 2585 12905 2619
rect 12939 2585 13001 2619
rect 13035 2585 13097 2619
rect 13131 2585 13193 2619
rect 13227 2585 13289 2619
rect 13323 2585 13385 2619
rect 13419 2585 13481 2619
rect 13515 2617 17682 2619
rect 13515 2585 13923 2617
rect 5634 2583 13923 2585
rect 13957 2583 14019 2617
rect 14053 2583 14115 2617
rect 14149 2583 14211 2617
rect 14245 2583 14307 2617
rect 14341 2583 14403 2617
rect 14437 2583 14499 2617
rect 14533 2583 14595 2617
rect 14629 2583 14691 2617
rect 14725 2583 14787 2617
rect 14821 2583 14883 2617
rect 14917 2583 14979 2617
rect 15013 2583 15075 2617
rect 15109 2583 15171 2617
rect 15205 2583 15267 2617
rect 15301 2583 15363 2617
rect 15397 2583 15459 2617
rect 15493 2583 15555 2617
rect 15589 2613 17682 2617
rect 15589 2583 15985 2613
rect 5634 2579 15985 2583
rect 16019 2579 16081 2613
rect 16115 2579 16177 2613
rect 16211 2579 16273 2613
rect 16307 2579 16369 2613
rect 16403 2579 16465 2613
rect 16499 2579 16561 2613
rect 16595 2579 16657 2613
rect 16691 2579 16753 2613
rect 16787 2579 16849 2613
rect 16883 2579 16945 2613
rect 16979 2579 17041 2613
rect 17075 2579 17137 2613
rect 17171 2579 17233 2613
rect 17267 2579 17329 2613
rect 17363 2579 17425 2613
rect 17459 2579 17521 2613
rect 17555 2579 17617 2613
rect 17651 2579 17682 2613
rect 5634 2578 17682 2579
rect 5634 2565 7362 2578
rect 7696 2561 9424 2578
rect 9756 2574 15620 2578
rect 9756 2557 11484 2574
rect 11818 2553 13546 2574
rect 13892 2551 15620 2574
rect 15954 2547 17682 2578
rect 22544 2616 22820 2634
rect 22544 2603 22658 2616
rect 22712 2603 22820 2616
rect 22544 2569 22573 2603
rect 22607 2569 22658 2603
rect 22712 2569 22757 2603
rect 22791 2569 22820 2603
rect 22544 2556 22658 2569
rect 22712 2556 22820 2569
rect 22544 2538 22820 2556
rect 23168 2604 23444 2632
rect 23168 2601 23284 2604
rect 23342 2601 23444 2604
rect 23168 2567 23197 2601
rect 23231 2567 23284 2601
rect 23342 2567 23381 2601
rect 23415 2567 23444 2601
rect 23168 2550 23284 2567
rect 23342 2550 23444 2567
rect 23168 2536 23444 2550
rect 23776 2589 24236 2620
rect 23776 2555 23805 2589
rect 23839 2555 23897 2589
rect 23931 2588 23989 2589
rect 24023 2588 24081 2589
rect 23931 2555 23980 2588
rect 24042 2555 24081 2588
rect 24115 2555 24173 2589
rect 24207 2555 24236 2589
rect 23776 2532 23980 2555
rect 24042 2532 24236 2555
rect 23776 2524 24236 2532
rect 24600 2594 25244 2606
rect 24600 2575 24892 2594
rect 24954 2575 25244 2594
rect 24600 2541 24629 2575
rect 24663 2541 24721 2575
rect 24755 2541 24813 2575
rect 24847 2541 24892 2575
rect 24954 2541 24997 2575
rect 25031 2541 25089 2575
rect 25123 2541 25181 2575
rect 25215 2541 25244 2575
rect 24600 2538 24892 2541
rect 24954 2538 25244 2541
rect 24600 2510 25244 2538
rect 30392 174 30508 2758
rect 30390 144 30514 174
rect 30390 68 30408 144
rect 30482 68 30514 144
rect 30390 34 30514 68
<< via1 >>
rect 904 4420 958 4486
rect 8192 4138 8244 4142
rect 8192 4096 8220 4138
rect 8220 4096 8244 4138
rect 8192 4090 8244 4096
rect 344 3740 438 3830
rect 366 3228 442 3320
rect 2132 2936 2184 2988
rect 1000 2582 1066 2660
rect 22654 3147 22706 3158
rect 22654 3113 22665 3147
rect 22665 3113 22699 3147
rect 22699 3113 22706 3147
rect 22654 3106 22706 3113
rect 23268 3145 23326 3152
rect 23268 3111 23289 3145
rect 23289 3111 23323 3145
rect 23323 3111 23326 3145
rect 23268 3096 23326 3111
rect 23982 3133 24040 3152
rect 23982 3099 23989 3133
rect 23989 3099 24023 3133
rect 24023 3099 24040 3133
rect 23982 3096 24040 3099
rect 24914 3119 24972 3138
rect 24914 3085 24939 3119
rect 24939 3085 24972 3119
rect 24914 3082 24972 3085
rect 22658 2603 22712 2616
rect 22658 2569 22665 2603
rect 22665 2569 22699 2603
rect 22699 2569 22712 2603
rect 22658 2556 22712 2569
rect 23284 2601 23342 2604
rect 23284 2567 23289 2601
rect 23289 2567 23323 2601
rect 23323 2567 23342 2601
rect 23284 2550 23342 2567
rect 23980 2555 23989 2588
rect 23989 2555 24023 2588
rect 24023 2555 24042 2588
rect 23980 2532 24042 2555
rect 24892 2575 24954 2594
rect 24892 2541 24905 2575
rect 24905 2541 24939 2575
rect 24939 2541 24954 2575
rect 24892 2538 24954 2541
rect 30408 68 30482 144
<< metal2 >>
rect 890 4486 972 4516
rect 890 4420 904 4486
rect 960 4420 972 4486
rect 890 4386 972 4420
rect 2126 4142 8254 4174
rect 2126 4090 8192 4142
rect 8244 4090 8254 4142
rect 2126 4070 8254 4090
rect 2126 4044 2244 4070
rect 294 3830 484 3880
rect 294 3740 344 3830
rect 438 3740 484 3830
rect 294 3684 484 3740
rect 354 3320 466 3390
rect 354 3228 366 3320
rect 442 3228 466 3320
rect 354 3166 466 3228
rect 2128 2994 2188 4044
rect 22580 3162 22786 3168
rect 22580 3106 22654 3162
rect 22712 3106 22786 3162
rect 22580 3082 22786 3106
rect 23192 3152 23398 3172
rect 23192 3096 23268 3152
rect 23326 3096 23398 3152
rect 23192 3086 23398 3096
rect 23908 3152 24114 3168
rect 23908 3096 23982 3152
rect 24040 3096 24114 3152
rect 23908 3082 24114 3096
rect 24848 3138 25054 3150
rect 24848 3082 24914 3138
rect 24972 3082 25054 3138
rect 24848 3064 25054 3082
rect 2104 2988 2194 2994
rect 2104 2936 2132 2988
rect 2184 2936 2194 2988
rect 2104 2922 2194 2936
rect 966 2660 1096 2704
rect 966 2582 1000 2660
rect 1066 2582 1096 2660
rect 966 2522 1096 2582
rect 22546 2616 22794 2630
rect 22546 2556 22658 2616
rect 22714 2556 22794 2616
rect 22546 2534 22794 2556
rect 23178 2606 23426 2628
rect 23178 2550 23284 2606
rect 23342 2550 23426 2606
rect 23178 2532 23426 2550
rect 23870 2588 24118 2628
rect 23870 2532 23980 2588
rect 24042 2532 24118 2588
rect 24814 2594 25062 2600
rect 24814 2538 24892 2594
rect 24954 2538 25062 2594
rect 24814 2504 25062 2538
rect 30390 144 30514 174
rect 30390 68 30408 144
rect 30482 68 30514 144
rect 30390 34 30514 68
<< via2 >>
rect 904 4420 958 4486
rect 958 4420 960 4486
rect 344 3740 438 3830
rect 366 3228 442 3320
rect 22654 3158 22712 3162
rect 22654 3106 22706 3158
rect 22706 3106 22712 3158
rect 23268 3096 23326 3152
rect 23982 3096 24040 3152
rect 24914 3082 24972 3138
rect 1000 2582 1066 2660
rect 22658 2556 22712 2616
rect 22712 2556 22714 2616
rect 23284 2604 23342 2606
rect 23284 2550 23342 2604
rect 23980 2532 24042 2588
rect 24892 2538 24954 2594
rect 30408 68 30482 144
<< metal3 >>
rect 890 4486 972 4516
rect 890 4420 904 4486
rect 968 4420 972 4486
rect 890 4386 972 4420
rect 294 3830 484 3880
rect 294 3740 344 3830
rect 438 3740 484 3830
rect 294 3684 484 3740
rect 464 3566 25256 3608
rect 464 3500 508 3566
rect 572 3500 25256 3566
rect 464 3450 25256 3500
rect 524 3406 25256 3450
rect 354 3320 466 3390
rect 354 3228 366 3320
rect 442 3228 466 3320
rect 354 3166 466 3228
rect 22591 3162 22793 3406
rect 22591 3106 22654 3162
rect 22712 3106 22793 3162
rect 22591 3085 22793 3106
rect 23181 3152 23383 3406
rect 23181 3096 23268 3152
rect 23326 3096 23383 3152
rect 23181 3077 23383 3096
rect 23915 3152 24117 3406
rect 23915 3096 23982 3152
rect 24040 3096 24117 3152
rect 23915 3069 24117 3096
rect 24841 3138 25043 3406
rect 24841 3082 24914 3138
rect 24972 3082 25043 3138
rect 24841 3055 25043 3082
rect 966 2660 1096 2704
rect 966 2582 1000 2660
rect 1066 2582 1096 2660
rect 966 2522 1096 2582
rect 22493 2616 22791 2627
rect 22493 2556 22658 2616
rect 22714 2556 22791 2616
rect 22493 2266 22791 2556
rect 23149 2606 23447 2625
rect 23149 2550 23284 2606
rect 23342 2550 23447 2606
rect 23149 2266 23447 2550
rect 23843 2588 24141 2613
rect 23843 2532 23980 2588
rect 24042 2532 24141 2588
rect 23843 2266 24141 2532
rect 24783 2594 25081 2603
rect 24783 2538 24892 2594
rect 24954 2538 25081 2594
rect 24783 2266 25081 2538
rect 1006 2154 25200 2266
rect 1006 2052 1048 2154
rect 1146 2052 25200 2154
rect 1006 1968 25200 2052
rect 30390 144 30514 174
rect 30390 68 30408 144
rect 30482 68 30514 144
rect 30390 34 30514 68
<< via3 >>
rect 904 4420 960 4486
rect 960 4420 968 4486
rect 344 3740 438 3830
rect 508 3500 572 3566
rect 366 3228 442 3320
rect 1000 2582 1066 2660
rect 1048 2052 1146 2154
rect 30408 68 30482 144
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 3830 600 44152
rect 200 3740 344 3830
rect 438 3740 600 3830
rect 200 3566 600 3740
rect 200 3500 508 3566
rect 572 3500 600 3566
rect 200 3320 600 3500
rect 200 3228 366 3320
rect 442 3228 600 3320
rect 200 1000 600 3228
rect 800 4486 1200 44152
rect 800 4420 904 4486
rect 968 4420 1200 4486
rect 800 2660 1200 4420
rect 800 2582 1000 2660
rect 1066 2582 1200 2660
rect 800 2154 1200 2582
rect 800 2052 1048 2154
rect 1146 2052 1200 2154
rect 800 1000 1200 2052
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 144 30542 200
rect 30362 68 30408 144
rect 30482 68 30542 144
rect 30362 0 30542 68
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel comment s 3560 2616 3560 2616 4 fa_1
flabel pwell s 3560 2616 5288 2665 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 3560 3233 5288 3282 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 3560 3233 5288 3282 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 3560 2616 5288 2665 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 4455 2858 4489 2892 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 4935 2932 4969 2966 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 3591 2710 3625 2744 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 3591 2784 3625 2818 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 1498 2620 1498 2620 4 fa_1
flabel pwell s 1498 2620 3226 2669 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 1498 3237 3226 3286 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 2297 2936 2331 2970 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel metal1 s 1498 3237 3226 3286 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 1498 2620 3226 2669 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2393 2862 2427 2896 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2873 2936 2907 2970 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1529 2714 1563 2748 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1529 2788 1563 2822 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 5665 2782 5699 2816 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 5665 2708 5699 2742 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 7009 2930 7043 2964 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 6529 2856 6563 2890 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 5634 2614 7362 2663 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 5634 3231 7362 3280 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel nwell s 5634 3231 7362 3280 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 5634 2614 7362 2663 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 5634 2614 5634 2614 4 fa_1
flabel locali s 7727 2778 7761 2812 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 7727 2704 7761 2738 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 9071 2926 9105 2960 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 8591 2852 8625 2886 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 7696 2610 9424 2659 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 7696 3227 9424 3276 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel nwell s 7696 3227 9424 3276 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 7696 2610 9424 2659 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 7696 2610 7696 2610 4 fa_1
rlabel comment s 13892 2600 13892 2600 4 fa_1
flabel pwell s 13892 2600 15620 2649 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 13892 3217 15620 3266 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 13892 3217 15620 3266 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 13892 2600 15620 2649 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 14787 2842 14821 2876 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 15267 2916 15301 2950 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 13923 2694 13957 2728 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 13923 2768 13957 2802 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 15954 2596 15954 2596 4 fa_1
flabel pwell s 15954 2596 17682 2645 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 15954 3213 17682 3262 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 15954 3213 17682 3262 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 15954 2596 17682 2645 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 16849 2838 16883 2872 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 17329 2912 17363 2946 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 17617 2690 17651 2724 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2764 17651 2798 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2838 17651 2872 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2912 17651 2946 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 2986 17651 3020 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 3060 17651 3094 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 17617 3134 17651 3168 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 15985 2690 16019 2724 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 15985 2764 16019 2798 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 11818 2602 11818 2602 4 fa_1
flabel pwell s 11818 2602 13546 2651 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 11818 3219 13546 3268 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 11818 3219 13546 3268 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 11818 2602 13546 2651 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 12713 2844 12747 2878 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 13193 2918 13227 2952 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 11849 2696 11883 2730 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 11849 2770 11883 2804 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment s 9756 2606 9756 2606 4 fa_1
flabel pwell s 9756 2606 11484 2655 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 9756 3223 11484 3272 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 9756 3223 11484 3272 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 9756 2606 11484 2655 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 10651 2848 10685 2882 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 11131 2922 11165 2956 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 9787 2700 9821 2734 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 9787 2774 9821 2808 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
rlabel comment 1498 2620 1498 2620 4 sky130_fd_sc_hs__fa_1_0.fa_1
flabel pwell 1498 2620 3226 2669 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_0.VNB
flabel nwell 1498 3237 3226 3286 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_0.VPB
flabel metal1 2297 2936 2331 2970 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.CIN
flabel metal1 1498 3237 3226 3286 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.VPWR
flabel metal1 1498 2620 3226 2669 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.VGND
flabel locali 2393 2862 2427 2896 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.A
flabel locali 2873 2936 2907 2970 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.B
flabel locali 3161 2714 3195 2748 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.COUT
flabel locali 3161 2788 3195 2822 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.COUT
flabel locali 3161 2862 3195 2896 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.COUT
flabel locali 3161 2936 3195 2970 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.COUT
flabel locali 3161 3010 3195 3044 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.COUT
flabel locali 3161 3084 3195 3118 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.COUT
flabel locali 3161 3158 3195 3192 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.COUT
flabel locali 1529 2714 1563 2748 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.SUM
flabel locali 1529 2788 1563 2822 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_0.SUM
rlabel comment 3560 2616 3560 2616 4 sky130_fd_sc_hs__fa_1_1.fa_1
flabel pwell 3560 2616 5288 2665 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_1.VNB
flabel nwell 3560 3233 5288 3282 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_1.VPB
flabel metal1 4359 2932 4393 2966 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.CIN
flabel metal1 3560 3233 5288 3282 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.VPWR
flabel metal1 3560 2616 5288 2665 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.VGND
flabel locali 4455 2858 4489 2892 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.A
flabel locali 4935 2932 4969 2966 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.B
flabel locali 5223 2710 5257 2744 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.COUT
flabel locali 5223 2784 5257 2818 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.COUT
flabel locali 5223 2858 5257 2892 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.COUT
flabel locali 5223 2932 5257 2966 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.COUT
flabel locali 5223 3006 5257 3040 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.COUT
flabel locali 5223 3080 5257 3114 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.COUT
flabel locali 5223 3154 5257 3188 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.COUT
flabel locali 3591 2710 3625 2744 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.SUM
flabel locali 3591 2784 3625 2818 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_1.SUM
rlabel comment 5634 2614 5634 2614 4 sky130_fd_sc_hs__fa_1_3.fa_1
flabel pwell 5634 2614 7362 2663 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_3.VNB
flabel nwell 5634 3231 7362 3280 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_3.VPB
flabel metal1 6433 2930 6467 2964 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.CIN
flabel metal1 5634 3231 7362 3280 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.VPWR
flabel metal1 5634 2614 7362 2663 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.VGND
flabel locali 6529 2856 6563 2890 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.A
flabel locali 7009 2930 7043 2964 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.B
flabel locali 7297 2708 7331 2742 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.COUT
flabel locali 7297 2782 7331 2816 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.COUT
flabel locali 7297 2856 7331 2890 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.COUT
flabel locali 7297 2930 7331 2964 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.COUT
flabel locali 7297 3004 7331 3038 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.COUT
flabel locali 7297 3078 7331 3112 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.COUT
flabel locali 7297 3152 7331 3186 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.COUT
flabel locali 5665 2708 5699 2742 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.SUM
flabel locali 5665 2782 5699 2816 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_3.SUM
rlabel comment 7696 2610 7696 2610 4 sky130_fd_sc_hs__fa_1_2.fa_1
flabel pwell 7696 2610 9424 2659 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_2.VNB
flabel nwell 7696 3227 9424 3276 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_2.VPB
flabel metal1 8495 2926 8529 2960 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.CIN
flabel metal1 7696 3227 9424 3276 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.VPWR
flabel metal1 7696 2610 9424 2659 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.VGND
flabel locali 8591 2852 8625 2886 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.A
flabel locali 9071 2926 9105 2960 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.B
flabel locali 9359 2704 9393 2738 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.COUT
flabel locali 9359 2778 9393 2812 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.COUT
flabel locali 9359 2852 9393 2886 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.COUT
flabel locali 9359 2926 9393 2960 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.COUT
flabel locali 9359 3000 9393 3034 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.COUT
flabel locali 9359 3074 9393 3108 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.COUT
flabel locali 9359 3148 9393 3182 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.COUT
flabel locali 7727 2704 7761 2738 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.SUM
flabel locali 7727 2778 7761 2812 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_2.SUM
rlabel comment 8386 4452 8386 4452 8 sky130_fd_sc_hs__inv_2_0.inv_2
flabel pwell 8098 4403 8386 4452 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__inv_2_0.VNB
flabel nwell 8098 3786 8386 3835 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__inv_2_0.VPB
flabel metal1 8098 3786 8386 3835 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.VPWR
flabel metal1 8098 4403 8386 4452 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.VGND
flabel locali 8321 4102 8355 4136 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.A
flabel locali 8225 4324 8259 4358 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.Y
flabel locali 8225 4250 8259 4284 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.Y
flabel locali 8225 4176 8259 4210 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.Y
flabel locali 8225 4102 8259 4136 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.Y
flabel locali 8225 4028 8259 4062 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.Y
flabel locali 8225 3954 8259 3988 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.Y
flabel locali 8225 3880 8259 3914 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__inv_2_0.Y
rlabel comment 9756 2606 9756 2606 4 sky130_fd_sc_hs__fa_1_7.fa_1
flabel pwell 9756 2606 11484 2655 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_7.VNB
flabel nwell 9756 3223 11484 3272 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_7.VPB
flabel metal1 10555 2922 10589 2956 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.CIN
flabel metal1 9756 3223 11484 3272 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.VPWR
flabel metal1 9756 2606 11484 2655 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.VGND
flabel locali 10651 2848 10685 2882 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.A
flabel locali 11131 2922 11165 2956 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.B
flabel locali 11419 2700 11453 2734 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.COUT
flabel locali 11419 2774 11453 2808 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.COUT
flabel locali 11419 2848 11453 2882 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.COUT
flabel locali 11419 2922 11453 2956 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.COUT
flabel locali 11419 2996 11453 3030 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.COUT
flabel locali 11419 3070 11453 3104 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.COUT
flabel locali 11419 3144 11453 3178 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.COUT
flabel locali 9787 2700 9821 2734 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.SUM
flabel locali 9787 2774 9821 2808 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_7.SUM
rlabel comment 11818 2602 11818 2602 4 sky130_fd_sc_hs__fa_1_6.fa_1
flabel pwell 11818 2602 13546 2651 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_6.VNB
flabel nwell 11818 3219 13546 3268 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_6.VPB
flabel metal1 12617 2918 12651 2952 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.CIN
flabel metal1 11818 3219 13546 3268 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.VPWR
flabel metal1 11818 2602 13546 2651 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.VGND
flabel locali 12713 2844 12747 2878 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.A
flabel locali 13193 2918 13227 2952 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.B
flabel locali 13481 2696 13515 2730 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.COUT
flabel locali 13481 2770 13515 2804 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.COUT
flabel locali 13481 2844 13515 2878 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.COUT
flabel locali 13481 2918 13515 2952 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.COUT
flabel locali 13481 2992 13515 3026 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.COUT
flabel locali 13481 3066 13515 3100 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.COUT
flabel locali 13481 3140 13515 3174 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.COUT
flabel locali 11849 2696 11883 2730 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.SUM
flabel locali 11849 2770 11883 2804 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_6.SUM
rlabel comment 13892 2600 13892 2600 4 sky130_fd_sc_hs__fa_1_4.fa_1
flabel pwell 13892 2600 15620 2649 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_4.VNB
flabel nwell 13892 3217 15620 3266 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_4.VPB
flabel metal1 14691 2916 14725 2950 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.CIN
flabel metal1 13892 3217 15620 3266 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.VPWR
flabel metal1 13892 2600 15620 2649 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.VGND
flabel locali 14787 2842 14821 2876 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.A
flabel locali 15267 2916 15301 2950 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.B
flabel locali 15555 2694 15589 2728 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.COUT
flabel locali 15555 2768 15589 2802 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.COUT
flabel locali 15555 2842 15589 2876 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.COUT
flabel locali 15555 2916 15589 2950 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.COUT
flabel locali 15555 2990 15589 3024 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.COUT
flabel locali 15555 3064 15589 3098 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.COUT
flabel locali 15555 3138 15589 3172 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.COUT
flabel locali 13923 2694 13957 2728 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.SUM
flabel locali 13923 2768 13957 2802 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_4.SUM
rlabel comment 15954 2596 15954 2596 4 sky130_fd_sc_hs__fa_1_5.fa_1
flabel pwell 15954 2596 17682 2645 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_5.VNB
flabel nwell 15954 3213 17682 3262 0 FreeSans 200 0 0 0 sky130_fd_sc_hs__fa_1_5.VPB
flabel metal1 16753 2912 16787 2946 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.CIN
flabel metal1 15954 3213 17682 3262 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.VPWR
flabel metal1 15954 2596 17682 2645 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.VGND
flabel locali 16849 2838 16883 2872 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.A
flabel locali 17329 2912 17363 2946 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.B
flabel locali 17617 2690 17651 2724 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.COUT
flabel locali 17617 2764 17651 2798 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.COUT
flabel locali 17617 2838 17651 2872 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.COUT
flabel locali 17617 2912 17651 2946 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.COUT
flabel locali 17617 2986 17651 3020 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.COUT
flabel locali 17617 3060 17651 3094 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.COUT
flabel locali 17617 3134 17651 3168 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.COUT
flabel locali 15985 2690 16019 2724 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.SUM
flabel locali 15985 2764 16019 2798 0 FreeSans 340 0 0 0 sky130_fd_sc_hs__fa_1_5.SUM
flabel locali 25173 2711 25207 2745 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.Y
flabel locali 25173 2779 25207 2813 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.Y
flabel locali 25173 2847 25207 2881 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.Y
flabel locali 24629 2779 24663 2813 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel locali 24897 2779 24931 2813 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel locali 24989 2779 25023 2813 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel locali 25081 2779 25115 2813 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel nwell 24629 3085 24663 3119 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VPB
flabel pwell 24629 2541 24663 2575 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VNB
flabel metal1 24629 3085 24663 3119 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VPWR
flabel metal1 24629 2541 24663 2575 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VGND
rlabel comment 24600 2558 24600 2558 4 sky130_fd_sc_hd__inv_6_0.inv_6
rlabel metal1 24600 2510 25244 2606 1 sky130_fd_sc_hd__inv_6_0.VGND
rlabel metal1 24600 3054 25244 3150 1 sky130_fd_sc_hd__inv_6_0.VPWR
flabel locali 24173 2725 24207 2759 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.Y
flabel locali 24173 2793 24207 2827 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.Y
flabel locali 24173 2861 24207 2895 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.Y
flabel locali 23805 2793 23839 2827 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel locali 23897 2793 23931 2827 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel locali 23989 2793 24023 2827 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel locali 24081 2793 24115 2827 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel nwell 23805 3099 23839 3133 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VPB
flabel pwell 23805 2555 23839 2589 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VNB
flabel metal1 23805 3099 23839 3133 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VPWR
flabel metal1 23805 2555 23839 2589 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VGND
rlabel comment 23776 2572 23776 2572 4 sky130_fd_sc_hd__inv_4_0.inv_4
rlabel metal1 23776 2524 24236 2620 1 sky130_fd_sc_hd__inv_4_0.VGND
rlabel metal1 23776 3068 24236 3164 1 sky130_fd_sc_hd__inv_4_0.VPWR
flabel locali 23197 2805 23231 2839 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.A
flabel locali 23289 2737 23323 2771 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.Y
flabel locali 23289 2873 23323 2907 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.Y
flabel locali 23289 2805 23323 2839 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.Y
flabel nwell 23197 3111 23231 3145 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VPB
flabel pwell 23197 2567 23231 2601 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VNB
flabel metal1 23197 3111 23231 3145 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VPWR
flabel metal1 23197 2567 23231 2601 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VGND
rlabel comment 23168 2584 23168 2584 4 sky130_fd_sc_hd__inv_2_0.inv_2
rlabel metal1 23168 2536 23444 2632 1 sky130_fd_sc_hd__inv_2_0.VGND
rlabel metal1 23168 3080 23444 3176 1 sky130_fd_sc_hd__inv_2_0.VPWR
flabel locali 22708 2875 22742 2909 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0.Y
flabel locali 22708 2807 22742 2841 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0.Y
flabel locali 22616 2807 22650 2841 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0.A
flabel nwell 22573 3113 22607 3147 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0.VPB
flabel pwell 22573 2569 22607 2603 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0.VNB
flabel metal1 22573 2569 22607 2603 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0.VGND
flabel metal1 22573 3113 22607 3147 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0.VPWR
rlabel comment 22544 2586 22544 2586 4 sky130_fd_sc_hd__inv_1_0.inv_1
rlabel metal1 22544 2538 22820 2634 1 sky130_fd_sc_hd__inv_1_0.VGND
rlabel metal1 22544 3082 22820 3178 1 sky130_fd_sc_hd__inv_1_0.VPWR
<< end >>
