* NGSPICE file created from tt_um_ohmy90_ringOscillator.ext - technology: sky130B

.subckt sky130_fd_sc_hs__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM a_1100_75# a_1107_347#
+ a_318_389# a_315_75# a_916_347# a_69_260# a_936_75# a_465_249# a_237_75# a_501_75#
+ a_509_347# a_217_368#
X0 a_465_249# B a_936_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=3584,184
X1 a_501_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=6763,255 d=3584,184
X2 a_318_389# B a_217_368# VPB sky130_fd_pr__pfet_01v8 ad=0.19588 pd=1.565 as=0.18669 ps=1.46 w=1 l=0.15
**devattr s=7467,292 d=7835,313
X3 VPWR CIN a_509_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.1725 ps=1.345 w=1 l=0.15
**devattr s=7100,271 d=6200,262
X4 a_69_260# CIN a_315_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=4992,206
X5 a_501_75# a_465_249# a_69_260# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.1248 ps=1.03 w=0.64 l=0.15
**devattr s=4992,206 d=4608,200
X6 VGND A a_1100_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.29627 ps=1.75667 w=0.64 l=0.15
**devattr s=14384,346 d=8491,282
X7 VGND a_69_260# SUM VNB sky130_fd_pr__nfet_01v8_lvt ad=0.20595 pd=1.54456 as=0.2109 ps=2.05 w=0.74 l=0.15
**devattr s=8436,410 d=7663,279
X8 VGND CIN a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.1024 ps=0.96 w=0.64 l=0.15
**devattr s=3584,184 d=6336,227
X9 a_237_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=7663,279 d=3072,176
X10 a_509_347# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=9745,328 d=7100,271
X11 COUT a_465_249# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.26955 ps=1.84485 w=1.12 l=0.15
**devattr s=13216,566 d=12768,562
X12 a_465_249# B a_916_347# VPB sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1775 ps=1.355 w=1 l=0.15
**devattr s=7100,271 d=6000,260
X13 a_1107_347# CIN a_465_249# VPB sky130_fd_pr__pfet_01v8 ad=0.26 pd=1.85333 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6000,260 d=8900,289
X14 VPWR A a_1107_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.26 ps=1.85333 w=1 l=0.15
**devattr s=8900,289 d=13962,352
X15 COUT a_465_249# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.20595 ps=1.54456 w=0.74 l=0.15
**devattr s=7844,402 d=7992,404
X16 a_1100_75# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.29627 pd=1.75667 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=8491,282 d=6784,362
X17 a_509_347# a_465_249# a_69_260# VPB sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6000,260 d=6700,267
X18 a_217_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.18669 pd=1.46 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=7960,297 d=7467,292
X19 a_916_347# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1775 pd=1.355 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=6200,262 d=7100,271
X20 a_936_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=6336,227 d=3072,176
X21 a_69_260# CIN a_318_389# VPB sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.19588 ps=1.565 w=1 l=0.15
**devattr s=7835,313 d=6000,260
X22 a_1100_75# CIN a_465_249# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.29627 pd=1.75667 as=0.0896 ps=0.92 w=0.64 l=0.15
**devattr s=3584,184 d=14384,346
X23 VPWR a_69_260# SUM VPB sky130_fd_pr__pfet_01v8 ad=0.26955 pd=1.84485 as=0.3192 ps=2.81 w=1.12 l=0.15
**devattr s=12768,562 d=7960,297
X24 VPWR B a_509_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.1725 ps=1.345 w=1 l=0.15
**devattr s=6700,267 d=9745,328
X25 a_1107_347# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.26 pd=1.85333 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=13962,352 d=13400,534
X26 a_315_75# B a_237_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=3072,176
X27 VGND B a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.1024 ps=0.96 w=0.64 l=0.15
**devattr s=4608,200 d=6763,255
C0 a_465_249# COUT 0.06928f
C1 CIN a_69_260# 0.10678f
C2 B a_69_260# 0.03966f
C3 VPB a_509_347# 0.00536f
C4 A a_315_75# 0.00252f
C5 a_465_249# a_501_75# 0.00555f
C6 a_1107_347# CIN 0.00192f
C7 CIN a_916_347# 0.0061f
C8 VGND CIN 0.13789f
C9 a_465_249# VPB 0.10732f
C10 a_1107_347# B 0.06557f
C11 VGND B 0.04033f
C12 SUM a_315_75# 0
C13 a_501_75# a_936_75# 0
C14 A a_217_368# 0
C15 VPWR a_69_260# 0.1278f
C16 a_1107_347# VPWR 0.21905f
C17 a_916_347# VPWR 0.01147f
C18 A SUM 0
C19 CIN B 0.19591f
C20 VGND VPWR 0.08465f
C21 a_1100_75# A 0.01955f
C22 a_1107_347# COUT 0
C23 CIN VPWR 0.13494f
C24 VGND COUT 0.07419f
C25 a_501_75# a_69_260# 0.02578f
C26 a_465_249# a_315_75# 0
C27 B VPWR 0.21956f
C28 VPB a_69_260# 0.04981f
C29 a_501_75# VGND 0.14715f
C30 a_1107_347# VPB 0.01475f
C31 VPB VGND 0.01302f
C32 A a_509_347# 0.01252f
C33 CIN COUT 0
C34 A a_465_249# 0.35643f
C35 B COUT 0.00688f
C36 A a_237_75# 0.00252f
C37 a_501_75# CIN 0.01116f
C38 A a_936_75# 0.00492f
C39 SUM a_237_75# 0
C40 VPB CIN 0.12323f
C41 a_501_75# B 0.00904f
C42 VPB B 0.62725f
C43 a_1100_75# a_465_249# 0.21113f
C44 VPWR COUT 0.12179f
C45 a_1100_75# a_936_75# 0
C46 a_315_75# a_69_260# 0.00702f
C47 VPB VPWR 0.24573f
C48 a_315_75# VGND 0.00207f
C49 a_217_368# a_69_260# 0.01644f
C50 a_465_249# a_509_347# 0.1366f
C51 A a_69_260# 0.27191f
C52 a_217_368# VGND 0.0017f
C53 a_465_249# a_237_75# 0
C54 A a_1107_347# 0.01477f
C55 A a_916_347# 0.0016f
C56 VPB COUT 0.01419f
C57 a_465_249# a_318_389# 0
C58 A VGND 0.13151f
C59 SUM a_69_260# 0.12447f
C60 a_315_75# CIN 0.00121f
C61 a_465_249# a_936_75# 0.00268f
C62 a_1100_75# a_69_260# 0
C63 SUM VGND 0.0376f
C64 a_1100_75# VGND 0.25139f
C65 A CIN 0.46738f
C66 A B 0.26846f
C67 SUM CIN 0
C68 SUM B 0
C69 a_509_347# a_69_260# 0.0624f
C70 a_1100_75# CIN 0.00368f
C71 a_217_368# VPWR 0.01541f
C72 a_1100_75# B 0.01175f
C73 a_465_249# a_69_260# 0.03228f
C74 A VPWR 0.04912f
C75 a_916_347# a_509_347# 0
C76 a_237_75# a_69_260# 0.00693f
C77 a_318_389# a_69_260# 0.02061f
C78 a_465_249# a_1107_347# 0.15034f
C79 a_465_249# a_916_347# 0.0195f
C80 a_465_249# VGND 0.12651f
C81 a_69_260# a_936_75# 0
C82 SUM VPWR 0.10504f
C83 VGND a_237_75# 0.00252f
C84 a_1100_75# VPWR 0.00321f
C85 VGND a_936_75# 0.0076f
C86 A COUT 0
C87 CIN a_509_347# 0.02394f
C88 B a_509_347# 0.02783f
C89 a_465_249# CIN 0.29824f
C90 a_465_249# B 0.27222f
C91 A a_501_75# 0.1337f
C92 CIN a_318_389# 0.00717f
C93 A VPB 0.14325f
C94 a_1100_75# COUT 0.00223f
C95 CIN a_936_75# 0.00177f
C96 SUM VPB 0.01283f
C97 VPWR a_509_347# 0.1543f
C98 a_465_249# VPWR 0.19408f
C99 VPWR a_237_75# 0
C100 VGND a_69_260# 0.15999f
C101 VPWR a_318_389# 0.01234f
C102 a_1107_347# VGND 0.00417f
C103 VGND VNB 0.99802f
C104 COUT VNB 0.11284f
C105 CIN VNB 0.31573f
C106 A VNB 0.49885f
C107 VPWR VNB 0.79012f
C108 SUM VNB 0.11694f
C109 B VNB 0.61239f
C110 VPB VNB 2.08861f
C111 a_1100_75# VNB 0.01137f
C112 a_501_75# VNB 0.00504f
C113 a_1107_347# VNB 0.00204f
C114 a_509_347# VNB 0.00129f
C115 a_465_249# VNB 0.30402f
C116 a_69_260# VNB 0.15472f
.ends

.subckt sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
**devattr s=8436,410 d=4144,204
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
**devattr s=6720,284 d=12768,562
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
**devattr s=4144,204 d=8436,410
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
**devattr s=12768,562 d=6720,284
C0 VPWR VPB 0.06315f
C1 Y A 0.11388f
C2 Y VGND 0.16424f
C3 A VGND 0.06173f
C4 VPWR Y 0.21165f
C5 VPB Y 0.00641f
C6 VPWR A 0.07533f
C7 VPB A 0.07759f
C8 VPWR VGND 0.0376f
C9 VPB VGND 0.00523f
C10 VGND VNB 0.30324f
C11 Y VNB 0.04146f
C12 VPWR VNB 0.26758f
C13 A VNB 0.30548f
C14 VPB VNB 0.40622f
.ends

.subckt tt_um_ohmy90_ringOscillator clk A B CIN ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
Xsky130_fd_sc_hs__fa_1_6 A B sky130_fd_sc_hs__fa_1_6/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_4/CIN
+ SUM a_12918_2677# a_12925_2949# a_12136_2991# a_12133_2677# a_12734_2949# a_11902_3194#
+ a_12754_2677# a_13432_3194# a_12055_2677# a_12319_2677# a_12327_2949# a_12035_2970#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_7 A B sky130_fd_sc_hs__fa_1_7/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_6/CIN
+ SUM a_10856_2681# a_10863_2953# a_10074_2995# a_10071_2681# a_10672_2953# a_9840_3198#
+ a_10692_2681# a_11370_3198# a_9993_2681# a_10257_2681# a_10265_2953# a_9973_2974#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_0 A B CIN A VNB VPB B sky130_fd_sc_hs__fa_1_1/CIN SUM a_2598_2695#
+ a_2605_2967# a_1816_3009# a_1813_2695# a_2414_2967# a_1582_3212# a_2434_2695# a_3112_3212#
+ a_1735_2695# a_1999_2695# a_2007_2967# a_1715_2988# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_1 A B sky130_fd_sc_hs__fa_1_1/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_3/CIN
+ SUM a_4660_2691# a_4667_2963# a_3878_3005# a_3875_2691# a_4476_2963# a_3644_3208#
+ a_4496_2691# a_5174_3208# a_3797_2691# a_4061_2691# a_4069_2963# a_3777_2984# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__inv_2_0 COUT A VNB sky130_fd_sc_hs__inv_2_0/VPB B CIN sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__fa_1_2 A B sky130_fd_sc_hs__fa_1_2/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_7/CIN
+ SUM a_8796_2685# a_8803_2957# a_8014_2999# a_8011_2685# a_8612_2957# a_7780_3202#
+ a_8632_2685# a_9310_3202# a_7933_2685# a_8197_2685# a_8205_2957# a_7913_2978# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_3 A B sky130_fd_sc_hs__fa_1_3/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_2/CIN
+ SUM a_6734_2689# a_6741_2961# a_5952_3003# a_5949_2689# a_6550_2961# a_5718_3206#
+ a_6570_2689# a_7248_3206# a_5871_2689# a_6135_2689# a_6143_2961# a_5851_2982# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_4 A B sky130_fd_sc_hs__fa_1_4/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_5/CIN
+ SUM a_14992_2675# a_14999_2947# a_14210_2989# a_14207_2675# a_14808_2947# a_13976_3192#
+ a_14828_2675# a_15506_3192# a_14129_2675# a_14393_2675# a_14401_2947# a_14109_2968#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_5 A B sky130_fd_sc_hs__fa_1_5/CIN A VNB VPB B COUT SUM a_17054_2671#
+ a_17061_2943# a_16272_2985# a_16269_2671# a_16870_2943# a_16038_3188# a_16890_2671#
+ a_17568_3188# a_16191_2671# a_16455_2671# a_16463_2943# a_16171_2964# sky130_fd_sc_hs__fa_1
C0 ui_in[1] ui_in[0] 0.03102f
C1 sky130_fd_sc_hs__fa_1_1/CIN SUM 0.07889f
C2 A a_16455_2671# 0.00604f
C3 a_5851_2982# B 0
C4 A a_16269_2671# 0
C5 uio_oe[0] uio_oe[1] 0.03102f
C6 B a_16870_2943# 0.00166f
C7 sky130_fd_sc_hs__fa_1_7/CIN a_9993_2681# 0.00127f
C8 B sky130_fd_sc_hs__fa_1_1/CIN 0.1412f
C9 sky130_fd_sc_hs__fa_1_3/CIN a_4660_2691# 0
C10 VPB a_5718_3206# 0
C11 a_7933_2685# sky130_fd_sc_hs__fa_1_2/CIN 0.00126f
C12 a_7780_3202# a_7248_3206# 0.00606f
C13 a_1715_2988# A 0
C14 B a_3797_2691# -0
C15 B a_4069_2963# 0.00165f
C16 B a_16463_2943# 0.00165f
C17 uio_out[5] uio_out[4] 0.03102f
C18 B a_4667_2963# 0.04723f
C19 uio_in[4] uio_in[3] 0.03102f
C20 CIN a_8014_2999# 0
C21 A a_2414_2967# 0
C22 B a_2598_2695# 0.00405f
C23 a_12319_2677# sky130_fd_sc_hs__fa_1_6/CIN 0
C24 sky130_fd_sc_hs__fa_1_6/CIN SUM 0.07889f
C25 a_1582_3212# A 0.00919f
C26 A a_12925_2949# -0.00169f
C27 VPB a_7248_3206# 0
C28 a_1715_2988# CIN 0.0017f
C29 a_9840_3198# VPB 0
C30 A COUT 0.041f
C31 a_12055_2677# sky130_fd_sc_hs__fa_1_6/CIN 0.00126f
C32 sky130_fd_sc_hs__fa_1_3/CIN a_6135_2689# 0
C33 A a_8205_2957# 0
C34 a_1582_3212# a_3112_3212# 0
C35 sky130_fd_sc_hs__fa_1_3/CIN sky130_fd_sc_hs__fa_1_2/CIN -0
C36 CIN a_2414_2967# 0.00304f
C37 A a_14828_2675# 0.003f
C38 B sky130_fd_sc_hs__fa_1_6/CIN 0.14229f
C39 a_9310_3202# SUM 0
C40 a_14129_2675# A 0
C41 uio_in[6] uio_in[5] 0.03102f
C42 B a_10074_2995# 0
C43 a_1582_3212# CIN 0.00855f
C44 A a_3875_2691# 0.00169f
C45 sky130_fd_sc_hs__fa_1_7/CIN a_11370_3198# 0
C46 sky130_fd_sc_hs__fa_1_7/CIN a_10672_2953# 0
C47 a_13976_3192# a_15506_3192# -0
C48 COUT CIN 0.07361f
C49 a_8205_2957# CIN 0
C50 B a_9310_3202# 0.02584f
C51 clk rst_n 0.03102f
C52 sky130_fd_sc_hs__fa_1_7/CIN a_8796_2685# -0
C53 a_11902_3194# sky130_fd_sc_hs__fa_1_6/CIN 0.06636f
C54 a_15506_3192# SUM 0
C55 a_9840_3198# a_10071_2681# 0
C56 a_4061_2691# A 0.06821f
C57 a_3875_2691# CIN 0
C58 B a_15506_3192# 0.0258f
C59 a_13976_3192# sky130_fd_sc_hs__fa_1_4/CIN 0.06234f
C60 sky130_fd_sc_hs__fa_1_5/CIN SUM 0.07889f
C61 sky130_fd_sc_hs__fa_1_7/CIN a_8803_2957# 0
C62 a_4061_2691# CIN 0
C63 a_7913_2978# sky130_fd_sc_hs__fa_1_2/CIN 0.00449f
C64 A a_14393_2675# 0.00604f
C65 SUM sky130_fd_sc_hs__fa_1_4/CIN 0.07548f
C66 a_8796_2685# sky130_fd_sc_hs__fa_1_2/CIN 0
C67 a_5174_3208# sky130_fd_sc_hs__fa_1_3/CIN 0.00595f
C68 uio_oe[3] uio_oe[4] 0.03102f
C69 B sky130_fd_sc_hs__fa_1_5/CIN 0.14093f
C70 A a_3112_3212# 0.01445f
C71 B sky130_fd_sc_hs__fa_1_4/CIN 0.1494f
C72 sky130_fd_sc_hs__fa_1_2/CIN a_8197_2685# 0
C73 B a_7933_2685# -0
C74 sky130_fd_sc_hs__fa_1_2/CIN a_8803_2957# -0
C75 A CIN 0.19782f
C76 A a_12327_2949# 0
C77 A a_6734_2689# 0.00618f
C78 sky130_fd_sc_hs__fa_1_3/CIN SUM 0.07548f
C79 B a_9993_2681# -0
C80 uo_out[7] uo_out[6] 0.03102f
C81 A a_5949_2689# 0
C82 CIN a_3112_3212# 0.03236f
C83 uio_out[1] uio_out[2] 0.03102f
C84 uo_out[3] uo_out[4] 0.03102f
C85 a_4476_2963# CIN 0
C86 B a_14808_2947# 0.00162f
C87 a_6734_2689# CIN 0
C88 B sky130_fd_sc_hs__fa_1_3/CIN 0.15023f
C89 sky130_fd_sc_hs__fa_1_6/CIN a_10856_2681# -0
C90 a_5949_2689# CIN 0
C91 a_16272_2985# sky130_fd_sc_hs__fa_1_5/CIN 0
C92 a_9840_3198# a_9310_3202# 0.00608f
C93 a_9310_3202# a_10856_2681# 0
C94 a_11370_3198# SUM 0
C95 a_10257_2681# a_11370_3198# 0
C96 a_14109_2968# sky130_fd_sc_hs__fa_1_4/CIN 0.0045f
C97 a_6741_2961# sky130_fd_sc_hs__fa_1_3/CIN 0
C98 B a_6143_2961# 0.00155f
C99 B a_10672_2953# 0.00166f
C100 B a_11370_3198# 0.02586f
C101 sky130_fd_sc_hs__fa_1_2/CIN a_8014_2999# 0
C102 A a_16171_2964# -0.0017f
C103 a_16038_3188# a_17568_3188# 0
C104 uio_out[6] uio_out[5] 0.03102f
C105 B a_7913_2978# 0
C106 B a_8796_2685# 0.00405f
C107 B a_16191_2671# -0
C108 a_11370_3198# a_11902_3194# 0.00606f
C109 B a_8197_2685# 0
C110 sky130_fd_sc_hs__fa_1_3/CIN a_5718_3206# 0.06234f
C111 B a_3777_2984# 0
C112 B a_8803_2957# 0.04723f
C113 a_8205_2957# sky130_fd_sc_hs__fa_1_2/CIN 0
C114 ui_in[1] ui_in[2] 0.03102f
C115 A a_10863_2953# -0.00169f
C116 B a_17061_2943# 0.04723f
C117 B a_2605_2967# 0.04723f
C118 sky130_fd_sc_hs__fa_1_3/CIN a_7248_3206# 0
C119 A a_4660_2691# 0.00617f
C120 uio_in[1] uio_in[2] 0.03102f
C121 sky130_fd_sc_hs__fa_1_3/CIN a_6550_2961# 0
C122 a_12133_2677# sky130_fd_sc_hs__fa_1_6/CIN 0
C123 a_14999_2947# A -0.00169f
C124 A a_14401_2947# 0
C125 a_4660_2691# a_3112_3212# 0
C126 sky130_fd_sc_hs__fa_1_7/CIN A 0.16537f
C127 B a_17054_2671# 0.00405f
C128 sky130_fd_sc_hs__fa_1_3/CIN a_5952_3003# 0
C129 VPB a_17568_3188# -0
C130 sky130_fd_sc_hs__fa_1_2/CIN a_8612_2957# 0
C131 a_16038_3188# VPB 0
C132 a_4660_2691# CIN 0
C133 B a_14992_2675# 0.00405f
C134 a_2007_2967# A 0.00166f
C135 uio_oe[5] uio_oe[4] 0.03102f
C136 B a_16455_2671# 0
C137 a_6143_2961# a_7248_3206# -0
C138 clk ena 0.03102f
C139 a_2007_2967# a_3112_3212# -0
C140 A a_6135_2689# 0.00604f
C141 A sky130_fd_sc_hs__fa_1_2/CIN 0.1614f
C142 a_9840_3198# a_11370_3198# -0
C143 a_2007_2967# CIN 0.01499f
C144 B a_8014_2999# 0
C145 a_8796_2685# a_7248_3206# 0
C146 a_11370_3198# a_10856_2681# -0
C147 B a_1715_2988# 0
C148 a_13976_3192# COUT 0
C149 A a_3644_3208# 0.05249f
C150 a_6135_2689# CIN 0
C151 a_6570_2689# a_7248_3206# 0
C152 a_1582_3212# SUM 0
C153 sky130_fd_sc_hs__fa_1_2/CIN CIN 0.00209f
C154 VPB a_7780_3202# 0
C155 sky130_fd_sc_hs__fa_1_2/CIN a_6734_2689# -0
C156 uio_out[2] uio_out[3] 0.03102f
C157 a_14129_2675# a_13976_3192# -0
C158 B a_2414_2967# 0.00148f
C159 a_5174_3208# a_4061_2691# 0
C160 a_3644_3208# a_3112_3212# 0.00606f
C161 a_17568_3188# a_16870_2943# 0
C162 A a_12734_2949# 0
C163 uio_in[7] uo_out[0] 0.03102f
C164 B a_1582_3212# 0.00152f
C165 B a_12925_2949# 0.04723f
C166 a_12918_2677# a_13432_3194# -0
C167 uo_out[3] uo_out[2] 0.03102f
C168 a_3644_3208# CIN 0.00209f
C169 B COUT 0.63711f
C170 B a_8205_2957# 0.00165f
C171 a_4496_2691# sky130_fd_sc_hs__fa_1_1/CIN -0
C172 a_16463_2943# a_17568_3188# -0
C173 B a_14129_2675# -0
C174 a_5174_3208# A 0.01477f
C175 a_13432_3194# VPB 0
C176 a_11902_3194# COUT 0
C177 a_2434_2695# a_1582_3212# -0
C178 a_13976_3192# a_14393_2675# 0
C179 B a_4061_2691# 0
C180 a_5174_3208# a_4476_2963# -0
C181 A a_13976_3192# -0
C182 a_5174_3208# CIN 0.00351f
C183 B a_8612_2957# 0.00166f
C184 a_5871_2689# sky130_fd_sc_hs__fa_1_3/CIN 0.00124f
C185 a_5174_3208# a_6734_2689# 0
C186 uio_in[6] uio_in[7] 0.03102f
C187 a_3878_3005# sky130_fd_sc_hs__fa_1_1/CIN 0
C188 A a_12319_2677# 0.00604f
C189 A SUM -0
C190 a_10257_2681# A 0.00604f
C191 a_12035_2970# sky130_fd_sc_hs__fa_1_6/CIN 0.00449f
C192 A a_12055_2677# 0
C193 a_3112_3212# SUM 0
C194 B a_14393_2675# 0
C195 B A 13.52898f
C196 VPB sky130_fd_sc_hs__fa_1_1/CIN 0.01675f
C197 sky130_fd_sc_hs__fa_1_7/CIN a_10863_2953# -0
C198 CIN SUM 0.0047f
C199 B a_3112_3212# 0.02517f
C200 B a_4476_2963# 0.00166f
C201 A a_11902_3194# -0
C202 a_16038_3188# a_15506_3192# 0.00606f
C203 B CIN 0.27871f
C204 uo_out[5] uo_out[4] 0.03102f
C205 a_1582_3212# a_1813_2695# 0
C206 B a_12327_2949# 0.00165f
C207 B a_6734_2689# 0.00405f
C208 a_12918_2677# sky130_fd_sc_hs__fa_1_6/CIN 0
C209 a_6741_2961# A -0.00169f
C210 a_2434_2695# A 0.00326f
C211 a_9840_3198# COUT 0
C212 a_17568_3188# sky130_fd_sc_hs__fa_1_5/CIN 0
C213 a_16038_3188# sky130_fd_sc_hs__fa_1_5/CIN 0.06636f
C214 a_9310_3202# a_7780_3202# 0
C215 a_2434_2695# a_3112_3212# 0
C216 a_14207_2675# sky130_fd_sc_hs__fa_1_4/CIN 0
C217 VPB sky130_fd_sc_hs__fa_1_6/CIN 0.01661f
C218 a_6741_2961# CIN 0.00105f
C219 a_1999_2695# a_1582_3212# 0
C220 sky130_fd_sc_hs__fa_1_7/CIN sky130_fd_sc_hs__fa_1_2/CIN -0
C221 a_2434_2695# CIN -0
C222 A a_14109_2968# -0.0017f
C223 a_13432_3194# sky130_fd_sc_hs__fa_1_6/CIN 0
C224 VPB a_9310_3202# 0
C225 A a_5718_3206# -0
C226 a_3797_2691# sky130_fd_sc_hs__fa_1_1/CIN 0.00126f
C227 a_4069_2963# sky130_fd_sc_hs__fa_1_1/CIN 0
C228 uio_oe[3] uio_oe[2] 0.03102f
C229 a_4667_2963# sky130_fd_sc_hs__fa_1_1/CIN -0
C230 uio_out[6] uio_out[7] 0.03102f
C231 A a_1813_2695# 0
C232 VPB a_15506_3192# 0
C233 a_2598_2695# sky130_fd_sc_hs__fa_1_1/CIN -0
C234 B a_16171_2964# 0
C235 a_5718_3206# CIN 0.00192f
C236 A a_7248_3206# 0.01078f
C237 a_5174_3208# a_4660_2691# -0
C238 a_11370_3198# a_10265_2953# -0
C239 a_9840_3198# A -0
C240 a_1813_2695# a_3112_3212# -0
C241 a_5718_3206# a_5949_2689# 0
C242 A a_10856_2681# 0.00618f
C243 sky130_fd_sc_hs__inv_2_0/VPB COUT 0.00689f
C244 uio_out[0] uo_out[7] 0.03102f
C245 VPB sky130_fd_sc_hs__fa_1_5/CIN 0.02401f
C246 VPB sky130_fd_sc_hs__fa_1_4/CIN 0.01809f
C247 uio_in[4] uio_in[5] 0.03102f
C248 CIN a_7248_3206# 0.0035f
C249 a_6734_2689# a_7248_3206# -0
C250 a_14210_2989# sky130_fd_sc_hs__fa_1_4/CIN 0
C251 a_1999_2695# A 0.00741f
C252 a_6550_2961# CIN 0
C253 a_13432_3194# sky130_fd_sc_hs__fa_1_4/CIN 0.00595f
C254 B a_12136_2991# 0
C255 a_1999_2695# a_3112_3212# -0
C256 uio_oe[2] uio_oe[1] 0.03102f
C257 a_5952_3003# CIN 0
C258 ui_in[3] ui_in[4] 0.03102f
C259 B a_10863_2953# 0.04723f
C260 sky130_fd_sc_hs__fa_1_7/CIN SUM 0.07963f
C261 a_1999_2695# CIN 0.00138f
C262 B a_4660_2691# 0.00405f
C263 sky130_fd_sc_hs__fa_1_7/CIN a_10257_2681# 0
C264 B a_14999_2947# 0.04723f
C265 VPB sky130_fd_sc_hs__fa_1_3/CIN 0.01799f
C266 uio_out[7] uio_oe[0] 0.03102f
C267 B a_14401_2947# 0.00155f
C268 ui_in[3] ui_in[2] 0.03102f
C269 sky130_fd_sc_hs__fa_1_7/CIN B 0.14154f
C270 a_5174_3208# a_3644_3208# 0
C271 sky130_fd_sc_hs__inv_2_0/VPB A 0
C272 a_12918_2677# a_11370_3198# 0
C273 B a_2007_2967# 0.00111f
C274 a_16870_2943# sky130_fd_sc_hs__fa_1_5/CIN 0
C275 sky130_fd_sc_hs__fa_1_2/CIN SUM 0.07889f
C276 B a_6135_2689# 0
C277 sky130_fd_sc_hs__inv_2_0/VPB CIN 0.0078f
C278 B sky130_fd_sc_hs__fa_1_2/CIN 0.14174f
C279 a_16463_2943# sky130_fd_sc_hs__fa_1_5/CIN 0
C280 a_3644_3208# SUM 0
C281 a_11370_3198# VPB 0.00733f
C282 a_17568_3188# a_16890_2671# -0
C283 a_5851_2982# sky130_fd_sc_hs__fa_1_3/CIN 0.0045f
C284 a_12133_2677# A 0
C285 uo_out[5] uo_out[6] 0.03102f
C286 B a_3644_3208# -0.00154f
C287 a_17568_3188# a_16455_2671# 0
C288 sky130_fd_sc_hs__fa_1_3/CIN sky130_fd_sc_hs__fa_1_1/CIN -0
C289 a_16269_2671# a_17568_3188# 0
C290 a_5871_2689# A 0
C291 B a_12734_2949# 0.00166f
C292 a_6741_2961# sky130_fd_sc_hs__fa_1_2/CIN 0
C293 sky130_fd_sc_hs__fa_1_6/CIN sky130_fd_sc_hs__fa_1_4/CIN -0
C294 sky130_fd_sc_hs__fa_1_6/CIN a_12754_2677# -0
C295 ui_in[5] ui_in[4] 0.03102f
C296 a_5174_3208# SUM 0
C297 a_4667_2963# sky130_fd_sc_hs__fa_1_3/CIN 0
C298 a_5871_2689# CIN 0
C299 a_5174_3208# B 0.02579f
C300 a_13976_3192# SUM 0
C301 a_5718_3206# a_6135_2689# 0
C302 sky130_fd_sc_hs__fa_1_7/CIN a_9840_3198# 0.06628f
C303 sky130_fd_sc_hs__fa_1_5/CIN a_15506_3192# 0.00578f
C304 a_17568_3188# COUT 0.02209f
C305 a_15506_3192# sky130_fd_sc_hs__fa_1_4/CIN 0
C306 ui_in[7] ui_in[6] 0.03102f
C307 sky130_fd_sc_hs__fa_1_7/CIN a_10856_2681# 0
C308 a_16038_3188# COUT 0
C309 B a_13976_3192# -0.00168f
C310 ui_in[7] uio_in[0] 0.03102f
C311 B a_12319_2677# 0
C312 B SUM -0
C313 a_10257_2681# B 0
C314 a_6135_2689# a_7248_3206# 0
C315 a_9973_2974# A -0.0017f
C316 sky130_fd_sc_hs__fa_1_2/CIN a_7248_3206# 0.00578f
C317 uo_out[1] uo_out[0] 0.03102f
C318 B a_12055_2677# -0
C319 sky130_fd_sc_hs__fa_1_5/CIN sky130_fd_sc_hs__fa_1_4/CIN -0
C320 a_3777_2984# sky130_fd_sc_hs__fa_1_1/CIN 0.00449f
C321 uio_oe[6] uio_oe[5] 0.03102f
C322 a_13432_3194# a_14992_2675# 0
C323 a_11902_3194# SUM 0
C324 A a_10265_2953# 0
C325 a_11370_3198# sky130_fd_sc_hs__fa_1_6/CIN 0.00642f
C326 a_1735_2695# a_1582_3212# -0
C327 a_2605_2967# sky130_fd_sc_hs__fa_1_1/CIN 0
C328 B a_11902_3194# -0.00159f
C329 a_5174_3208# a_5718_3206# 0.00609f
C330 A a_17568_3188# 0.01043f
C331 a_14808_2947# sky130_fd_sc_hs__fa_1_4/CIN 0
C332 uio_out[1] uio_out[0] 0.03102f
C333 a_6741_2961# B 0.04723f
C334 a_16038_3188# A -0
C335 a_14207_2675# A 0
C336 a_1582_3212# VPB 0
C337 a_8796_2685# a_9310_3202# -0
C338 a_12035_2970# A -0.0017f
C339 a_13976_3192# a_14109_2968# -0
C340 A a_8632_2685# 0.003f
C341 A a_4496_2691# 0.00346f
C342 VPB COUT 0.0186f
C343 B a_16272_2985# 0
C344 a_9310_3202# a_8197_2685# 0
C345 a_5718_3206# SUM 0
C346 a_13432_3194# COUT 0
C347 B a_14109_2968# 0
C348 a_4496_2691# CIN 0
C349 B a_5718_3206# -0.00163f
C350 a_12918_2677# A 0.00617f
C351 a_7248_3206# SUM 0
C352 a_1735_2695# A 0
C353 A a_7780_3202# -0
C354 a_9840_3198# SUM 0
C355 a_10257_2681# a_9840_3198# 0
C356 uio_in[1] uio_in[0] 0.03102f
C357 a_16191_2671# sky130_fd_sc_hs__fa_1_5/CIN 0.00126f
C358 a_1735_2695# a_3112_3212# 0
C359 B a_7248_3206# 0.02587f
C360 B a_9840_3198# -0.00151f
C361 a_3878_3005# CIN 0
C362 B a_6550_2961# 0.00162f
C363 sky130_fd_sc_hs__fa_1_3/CIN a_6143_2961# 0
C364 a_7780_3202# CIN 0.00188f
C365 A VPB -0.02614f
C366 B a_10856_2681# 0.00405f
C367 B a_5952_3003# 0
C368 VPB a_3112_3212# 0
C369 a_17061_2943# sky130_fd_sc_hs__fa_1_5/CIN -0
C370 a_17054_2671# a_15506_3192# 0
C371 a_13432_3194# A 0.01076f
C372 A a_1816_3009# 0
C373 B a_1999_2695# 0
C374 a_3875_2691# sky130_fd_sc_hs__fa_1_1/CIN 0
C375 VPB CIN 0.03018f
C376 a_14992_2675# a_15506_3192# -0
C377 sky130_fd_sc_hs__fa_1_3/CIN a_6570_2689# -0
C378 A a_10071_2681# 0
C379 a_4061_2691# sky130_fd_sc_hs__fa_1_1/CIN 0
C380 a_17054_2671# sky130_fd_sc_hs__fa_1_5/CIN 0
C381 a_1816_3009# CIN 0.00257f
C382 a_13432_3194# a_12327_2949# 0
C383 a_12925_2949# sky130_fd_sc_hs__fa_1_6/CIN -0
C384 sky130_fd_sc_hs__fa_1_5/CIN a_16890_2671# -0
C385 sky130_fd_sc_hs__fa_1_7/CIN a_9973_2974# 0.00447f
C386 a_5851_2982# A -0.0017f
C387 a_14992_2675# sky130_fd_sc_hs__fa_1_4/CIN 0
C388 uio_in[3] uio_in[2] 0.03102f
C389 sky130_fd_sc_hs__fa_1_5/CIN a_16455_2671# 0
C390 A sky130_fd_sc_hs__fa_1_1/CIN 0.16775f
C391 a_5718_3206# a_7248_3206# 0
C392 sky130_fd_sc_hs__inv_2_0/VPB B 0.01174f
C393 sky130_fd_sc_hs__fa_1_7/CIN a_10265_2953# 0
C394 a_16269_2671# sky130_fd_sc_hs__fa_1_5/CIN 0
C395 a_9310_3202# COUT 0
C396 a_9310_3202# a_8205_2957# 0
C397 a_5851_2982# CIN 0
C398 sky130_fd_sc_hs__fa_1_1/CIN a_3112_3212# 0.00578f
C399 a_3797_2691# A 0.00163f
C400 a_4069_2963# A 0
C401 a_16463_2943# A 0
C402 a_4476_2963# sky130_fd_sc_hs__fa_1_1/CIN 0
C403 a_4667_2963# A -0.00169f
C404 sky130_fd_sc_hs__fa_1_1/CIN CIN 0.00412f
C405 COUT a_15506_3192# 0
C406 A a_2598_2695# 0.00702f
C407 a_2598_2695# a_3112_3212# -0
C408 a_3797_2691# CIN 0
C409 a_4069_2963# CIN 0.00118f
C410 a_9310_3202# a_8612_2957# -0
C411 a_8011_2685# A 0
C412 a_4667_2963# CIN 0.00106f
C413 a_12925_2949# sky130_fd_sc_hs__fa_1_4/CIN 0
C414 A sky130_fd_sc_hs__fa_1_6/CIN 0.16195f
C415 COUT sky130_fd_sc_hs__fa_1_5/CIN 0
C416 a_2598_2695# CIN 0
C417 B a_5871_2689# -0
C418 a_14828_2675# sky130_fd_sc_hs__fa_1_4/CIN -0
C419 a_14129_2675# sky130_fd_sc_hs__fa_1_4/CIN 0.00124f
C420 a_10692_2681# A 0.003f
C421 A a_9310_3202# 0.01078f
C422 a_8011_2685# CIN 0
C423 a_8632_2685# sky130_fd_sc_hs__fa_1_2/CIN -0
C424 a_12327_2949# sky130_fd_sc_hs__fa_1_6/CIN 0
C425 a_15506_3192# a_14393_2675# 0
C426 A a_15506_3192# 0.01076f
C427 a_9310_3202# CIN 0
C428 sky130_fd_sc_hs__fa_1_7/CIN VPB 0.01694f
C429 uo_out[1] uo_out[2] 0.03102f
C430 sky130_fd_sc_hs__fa_1_2/CIN a_7780_3202# 0.06636f
C431 ui_in[5] ui_in[6] 0.03102f
C432 a_14393_2675# sky130_fd_sc_hs__fa_1_4/CIN 0
C433 A sky130_fd_sc_hs__fa_1_5/CIN 0.16338f
C434 A sky130_fd_sc_hs__fa_1_4/CIN 0.16183f
C435 a_7933_2685# A 0
C436 A a_12754_2677# 0.003f
C437 B a_9973_2974# 0
C438 a_5174_3208# a_4496_2691# -0
C439 a_5871_2689# a_5718_3206# -0
C440 VPB sky130_fd_sc_hs__fa_1_2/CIN 0.01668f
C441 sky130_fd_sc_hs__fa_1_7/CIN a_10071_2681# 0
C442 A a_9993_2681# 0
C443 a_11370_3198# COUT 0
C444 B a_10265_2953# 0.00166f
C445 a_7933_2685# CIN 0
C446 a_14207_2675# a_13976_3192# 0
C447 a_16038_3188# SUM 0
C448 a_4660_2691# sky130_fd_sc_hs__fa_1_1/CIN 0
C449 VPB a_3644_3208# 0
C450 A sky130_fd_sc_hs__fa_1_3/CIN 0.16269f
C451 B a_17568_3188# 0.02555f
C452 B a_16038_3188# -0.00159f
C453 B a_12035_2970# 0
C454 sky130_fd_sc_hs__fa_1_3/CIN CIN 0.00316f
C455 sky130_fd_sc_hs__fa_1_3/CIN a_6734_2689# 0
C456 a_13432_3194# a_12734_2949# 0
C457 sky130_fd_sc_hs__fa_1_6/CIN a_12136_2991# 0
C458 sky130_fd_sc_hs__fa_1_3/CIN a_5949_2689# 0
C459 A a_6143_2961# 0
C460 a_5174_3208# VPB 0
C461 sky130_fd_sc_hs__fa_1_6/CIN a_10863_2953# 0
C462 a_11370_3198# A 0.01078f
C463 a_7780_3202# SUM 0
C464 A a_7913_2978# -0.0017f
C465 a_8796_2685# A 0.00618f
C466 sky130_fd_sc_hs__fa_1_5/CIN a_16171_2964# 0.00449f
C467 a_17054_2671# COUT 0.00121f
C468 a_6143_2961# CIN 0.00118f
C469 B a_3878_3005# 0
C470 a_12918_2677# B 0.00405f
C471 VPB a_13976_3192# 0
C472 COUT a_16890_2671# 0
C473 B a_7780_3202# -0.00154f
C474 sky130_fd_sc_hs__fa_1_7/CIN sky130_fd_sc_hs__fa_1_6/CIN -0
C475 A a_16191_2671# 0
C476 a_3644_3208# sky130_fd_sc_hs__fa_1_1/CIN 0.06636f
C477 a_13976_3192# a_14210_2989# -0
C478 A a_6570_2689# 0.003f
C479 sky130_fd_sc_hs__fa_1_7/CIN a_10074_2995# 0
C480 A a_8197_2685# 0.00604f
C481 VPB SUM 0.01931f
C482 a_9840_3198# a_9973_2974# 0
C483 a_7913_2978# CIN 0
C484 sky130_fd_sc_hs__fa_1_7/CIN a_10692_2681# -0
C485 a_13432_3194# a_13976_3192# 0.00609f
C486 A a_3777_2984# -0.0017f
C487 uio_out[4] uio_out[3] 0.03102f
C488 sky130_fd_sc_hs__fa_1_7/CIN a_9310_3202# 0.00636f
C489 A a_8803_2957# -0.00169f
C490 a_13432_3194# a_12319_2677# 0
C491 a_13432_3194# SUM 0
C492 a_8011_2685# sky130_fd_sc_hs__fa_1_2/CIN 0
C493 B VPB 0.28716f
C494 B a_14210_2989# 0
C495 a_6570_2689# CIN 0
C496 A a_17061_2943# -0.00169f
C497 a_8197_2685# CIN 0
C498 uio_oe[6] uio_oe[7] 0.03102f
C499 a_2605_2967# A -0.00101f
C500 a_14401_2947# a_15506_3192# -0
C501 a_3777_2984# CIN 0
C502 a_5174_3208# sky130_fd_sc_hs__fa_1_1/CIN 0
C503 B a_1816_3009# 0
C504 B a_13432_3194# 0.02572f
C505 VPB a_11902_3194# 0
C506 a_9310_3202# sky130_fd_sc_hs__fa_1_2/CIN 0
C507 a_14999_2947# sky130_fd_sc_hs__fa_1_5/CIN 0
C508 a_17054_2671# A 0.00607f
C509 a_5174_3208# a_4069_2963# 0
C510 a_14999_2947# sky130_fd_sc_hs__fa_1_4/CIN 0
C511 a_2605_2967# CIN 0.00385f
C512 A a_16890_2671# 0.003f
C513 a_13432_3194# a_11902_3194# 0
C514 a_14992_2675# A 0.00618f
C515 a_14401_2947# sky130_fd_sc_hs__fa_1_4/CIN 0
C516 sky130_fd_sc_hs__fa_1_6/CIN a_12734_2949# 0
C517 rst_n ui_in[0] 0.03102f
C518 ua[1] VNB 0.1369f
C519 ua[2] VNB 0.1369f
C520 ua[3] VNB 0.1369f
C521 ua[4] VNB 0.1369f
C522 ua[5] VNB 0.1369f
C523 ua[6] VNB 0.1369f
C524 ua[7] VNB 0.1369f
C525 ena VNB 0.06503f
C526 clk VNB 0.03887f
C527 rst_n VNB 0.03887f
C528 ui_in[0] VNB 0.03887f
C529 ui_in[1] VNB 0.03887f
C530 ui_in[2] VNB 0.03887f
C531 ui_in[3] VNB 0.03887f
C532 ui_in[4] VNB 0.03887f
C533 ui_in[5] VNB 0.03887f
C534 ui_in[6] VNB 0.03887f
C535 ui_in[7] VNB 0.03887f
C536 uio_in[0] VNB 0.03887f
C537 uio_in[1] VNB 0.03887f
C538 uio_in[2] VNB 0.03887f
C539 uio_in[3] VNB 0.03887f
C540 uio_in[4] VNB 0.03887f
C541 uio_in[5] VNB 0.03887f
C542 uio_in[6] VNB 0.03887f
C543 uio_in[7] VNB 0.03887f
C544 uo_out[0] VNB 0.03887f
C545 uo_out[1] VNB 0.03887f
C546 uo_out[2] VNB 0.03887f
C547 uo_out[3] VNB 0.03887f
C548 uo_out[4] VNB 0.03887f
C549 uo_out[5] VNB 0.03887f
C550 uo_out[6] VNB 0.03887f
C551 uo_out[7] VNB 0.03887f
C552 uio_out[0] VNB 0.03887f
C553 uio_out[1] VNB 0.03887f
C554 uio_out[2] VNB 0.03887f
C555 uio_out[3] VNB 0.03887f
C556 uio_out[4] VNB 0.03887f
C557 uio_out[5] VNB 0.03887f
C558 uio_out[6] VNB 0.03887f
C559 uio_out[7] VNB 0.03887f
C560 uio_oe[0] VNB 0.03887f
C561 uio_oe[1] VNB 0.03887f
C562 uio_oe[2] VNB 0.03887f
C563 uio_oe[3] VNB 0.03887f
C564 uio_oe[4] VNB 0.03887f
C565 uio_oe[5] VNB 0.03887f
C566 uio_oe[6] VNB 0.03887f
C567 uio_oe[7] VNB 0.06503f
C568 a_17568_3188# VNB 0.30402f
C569 a_16038_3188# VNB 0.14774f
C570 a_15506_3192# VNB 0.2969f
C571 a_13976_3192# VNB 0.14781f
C572 a_13432_3194# VNB 0.29703f
C573 a_11902_3194# VNB 0.14774f
C574 a_11370_3198# VNB 0.27898f
C575 a_9840_3198# VNB 0.1477f
C576 a_9310_3202# VNB 0.29686f
C577 a_7780_3202# VNB 0.14774f
C578 a_7248_3206# VNB 0.2969f
C579 a_5718_3206# VNB 0.14781f
C580 B VNB 23.97779f
C581 a_5174_3208# VNB 0.29703f
C582 a_3644_3208# VNB 0.14774f
C583 a_3112_3212# VNB 0.2969f
C584 CIN VNB 2.25303f
C585 a_1582_3212# VNB 0.15472f
C586 COUT VNB 10.21649f
C587 a_17054_2671# VNB 0.01137f
C588 a_16455_2671# VNB 0.00504f
C589 a_17061_2943# VNB 0.00204f
C590 a_16463_2943# VNB 0.00129f
C591 sky130_fd_sc_hs__fa_1_5/CIN VNB 0.32654f
C592 a_14992_2675# VNB 0.01137f
C593 a_14393_2675# VNB 0.00504f
C594 a_14999_2947# VNB 0.00204f
C595 a_14401_2947# VNB 0.00129f
C596 sky130_fd_sc_hs__fa_1_2/CIN VNB 0.44151f
C597 sky130_fd_sc_hs__fa_1_3/CIN VNB 0.44533f
C598 a_6734_2689# VNB 0.01137f
C599 a_6135_2689# VNB 0.00504f
C600 a_6741_2961# VNB 0.00204f
C601 a_6143_2961# VNB 0.00129f
C602 a_8796_2685# VNB 0.01137f
C603 a_8197_2685# VNB 0.00504f
C604 a_8803_2957# VNB 0.00204f
C605 a_8205_2957# VNB 0.00129f
C606 sky130_fd_sc_hs__inv_2_0/VPB VNB 0.40622f
C607 a_4660_2691# VNB 0.01137f
C608 a_4061_2691# VNB 0.00504f
C609 a_4667_2963# VNB 0.00204f
C610 a_4069_2963# VNB 0.00129f
C611 sky130_fd_sc_hs__fa_1_1/CIN VNB 0.44129f
C612 A VNB 25.87713f
C613 SUM VNB 0.61793f
C614 VPB VNB 16.70885f
C615 a_2598_2695# VNB 0.01137f
C616 a_1999_2695# VNB 0.00504f
C617 a_2605_2967# VNB 0.00204f
C618 a_2007_2967# VNB 0.00129f
C619 sky130_fd_sc_hs__fa_1_6/CIN VNB 0.44099f
C620 sky130_fd_sc_hs__fa_1_7/CIN VNB 0.44071f
C621 a_10856_2681# VNB 0.01137f
C622 a_10257_2681# VNB 0.00504f
C623 a_10863_2953# VNB 0.00204f
C624 a_10265_2953# VNB 0.00129f
C625 sky130_fd_sc_hs__fa_1_4/CIN VNB 0.44615f
C626 a_12918_2677# VNB 0.01137f
C627 a_12319_2677# VNB 0.00504f
C628 a_12925_2949# VNB 0.00204f
C629 a_12327_2949# VNB 0.00129f
.ends

