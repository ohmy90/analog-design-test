* NGSPICE file created from tt_um_ohmy90_ringOscillator.ext - technology: sky130B

.subckt sky130_fd_sc_hs__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM a_1100_75# a_1107_347#
+ a_318_389# a_315_75# a_916_347# a_69_260# a_936_75# a_465_249# a_237_75# a_501_75#
+ a_509_347# a_217_368#
X0 a_465_249# B a_936_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=3584,184
X1 a_501_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=6763,255 d=3584,184
X2 a_318_389# B a_217_368# VPB sky130_fd_pr__pfet_01v8 ad=0.19588 pd=1.565 as=0.18669 ps=1.46 w=1 l=0.15
**devattr s=7467,292 d=7835,313
X3 VPWR CIN a_509_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.1725 ps=1.345 w=1 l=0.15
**devattr s=7100,271 d=6200,262
X4 a_69_260# CIN a_315_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=4992,206
X5 a_501_75# a_465_249# a_69_260# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1024 pd=0.96 as=0.1248 ps=1.03 w=0.64 l=0.15
**devattr s=4992,206 d=4608,200
X6 VGND A a_1100_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.29627 ps=1.75667 w=0.64 l=0.15
**devattr s=14384,346 d=8491,282
X7 VGND a_69_260# SUM VNB sky130_fd_pr__nfet_01v8_lvt ad=0.20595 pd=1.54456 as=0.2109 ps=2.05 w=0.74 l=0.15
**devattr s=8436,410 d=7663,279
X8 VGND CIN a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.1024 ps=0.96 w=0.64 l=0.15
**devattr s=3584,184 d=6336,227
X9 a_237_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=7663,279 d=3072,176
X10 a_509_347# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=9745,328 d=7100,271
X11 COUT a_465_249# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.26955 ps=1.84485 w=1.12 l=0.15
**devattr s=13216,566 d=12768,562
X12 a_465_249# B a_916_347# VPB sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1775 ps=1.355 w=1 l=0.15
**devattr s=7100,271 d=6000,260
X13 a_1107_347# CIN a_465_249# VPB sky130_fd_pr__pfet_01v8 ad=0.26 pd=1.85333 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6000,260 d=8900,289
X14 VPWR A a_1107_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.26 ps=1.85333 w=1 l=0.15
**devattr s=8900,289 d=13962,352
X15 COUT a_465_249# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.1998 pd=2.02 as=0.20595 ps=1.54456 w=0.74 l=0.15
**devattr s=7844,402 d=7992,404
X16 a_1100_75# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.29627 pd=1.75667 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=8491,282 d=6784,362
X17 a_509_347# a_465_249# a_69_260# VPB sky130_fd_pr__pfet_01v8 ad=0.1725 pd=1.345 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6000,260 d=6700,267
X18 a_217_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.18669 pd=1.46 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=7960,297 d=7467,292
X19 a_916_347# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.1775 pd=1.355 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=6200,262 d=7100,271
X20 a_936_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.17812 ps=1.33584 w=0.64 l=0.15
**devattr s=6336,227 d=3072,176
X21 a_69_260# CIN a_318_389# VPB sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.19588 ps=1.565 w=1 l=0.15
**devattr s=7835,313 d=6000,260
X22 a_1100_75# CIN a_465_249# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.29627 pd=1.75667 as=0.0896 ps=0.92 w=0.64 l=0.15
**devattr s=3584,184 d=14384,346
X23 VPWR a_69_260# SUM VPB sky130_fd_pr__pfet_01v8 ad=0.26955 pd=1.84485 as=0.3192 ps=2.81 w=1.12 l=0.15
**devattr s=12768,562 d=7960,297
X24 VPWR B a_509_347# VPB sky130_fd_pr__pfet_01v8 ad=0.24067 pd=1.64719 as=0.1725 ps=1.345 w=1 l=0.15
**devattr s=6700,267 d=9745,328
X25 a_1107_347# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0.26 pd=1.85333 as=0.24067 ps=1.64719 w=1 l=0.15
**devattr s=13962,352 d=13400,534
X26 a_315_75# B a_237_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.0768 pd=0.88 as=0.0768 ps=0.88 w=0.64 l=0.15
**devattr s=3072,176 d=3072,176
X27 VGND B a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt ad=0.17812 pd=1.33584 as=0.1024 ps=0.96 w=0.64 l=0.15
**devattr s=4608,200 d=6763,255
C0 A a_315_75# 0.00252f
C1 VGND A 0.13151f
C2 VPWR a_69_260# 0.1278f
C3 a_501_75# CIN 0.01116f
C4 a_916_347# CIN 0.0061f
C5 VPWR VPB 0.24573f
C6 a_1100_75# a_936_75# 0
C7 a_237_75# VPWR 0
C8 VGND a_1100_75# 0.25139f
C9 VGND VPWR 0.08465f
C10 B A 0.26846f
C11 a_1107_347# CIN 0.00192f
C12 a_465_249# COUT 0.06928f
C13 a_501_75# A 0.1337f
C14 a_465_249# a_509_347# 0.1366f
C15 a_916_347# A 0.0016f
C16 a_1100_75# B 0.01175f
C17 B VPWR 0.21956f
C18 VPB a_69_260# 0.04981f
C19 a_237_75# a_69_260# 0.00693f
C20 a_936_75# a_69_260# 0
C21 a_69_260# a_315_75# 0.00702f
C22 VGND a_69_260# 0.15999f
C23 a_1107_347# A 0.01477f
C24 a_916_347# VPWR 0.01147f
C25 VGND VPB 0.01302f
C26 a_465_249# CIN 0.29824f
C27 COUT CIN 0
C28 VGND a_237_75# 0.00252f
C29 VGND a_936_75# 0.0076f
C30 a_509_347# CIN 0.02394f
C31 VGND a_315_75# 0.00207f
C32 a_1107_347# VPWR 0.21905f
C33 B a_69_260# 0.03966f
C34 SUM CIN 0
C35 B VPB 0.62725f
C36 a_501_75# a_69_260# 0.02578f
C37 a_318_389# a_465_249# 0
C38 a_465_249# A 0.35643f
C39 VGND B 0.04033f
C40 A COUT 0
C41 a_509_347# A 0.01252f
C42 a_501_75# a_936_75# 0
C43 VGND a_501_75# 0.14715f
C44 a_465_249# a_1100_75# 0.21113f
C45 a_465_249# VPWR 0.19408f
C46 a_1100_75# COUT 0.00223f
C47 SUM A 0
C48 COUT VPWR 0.12179f
C49 a_1107_347# VPB 0.01475f
C50 a_509_347# VPWR 0.1543f
C51 a_318_389# CIN 0.00717f
C52 VGND a_1107_347# 0.00417f
C53 B a_501_75# 0.00904f
C54 A CIN 0.46738f
C55 a_217_368# A 0
C56 SUM VPWR 0.10504f
C57 a_1100_75# CIN 0.00368f
C58 a_465_249# a_69_260# 0.03228f
C59 VPWR CIN 0.13494f
C60 a_1107_347# B 0.06557f
C61 a_217_368# VPWR 0.01541f
C62 a_509_347# a_69_260# 0.0624f
C63 a_465_249# VPB 0.10732f
C64 COUT VPB 0.01419f
C65 a_509_347# VPB 0.00536f
C66 a_465_249# a_237_75# 0
C67 a_465_249# a_936_75# 0.00268f
C68 a_465_249# a_315_75# 0
C69 VGND a_465_249# 0.12651f
C70 SUM a_69_260# 0.12447f
C71 VGND COUT 0.07419f
C72 a_318_389# VPWR 0.01234f
C73 a_1100_75# A 0.01955f
C74 SUM VPB 0.01283f
C75 A VPWR 0.04912f
C76 SUM a_237_75# 0
C77 CIN a_69_260# 0.10678f
C78 a_217_368# a_69_260# 0.01644f
C79 SUM a_315_75# 0
C80 VGND SUM 0.0376f
C81 a_465_249# B 0.27222f
C82 CIN VPB 0.12323f
C83 B COUT 0.00688f
C84 a_509_347# B 0.02783f
C85 a_1100_75# VPWR 0.00321f
C86 a_936_75# CIN 0.00177f
C87 a_465_249# a_501_75# 0.00555f
C88 CIN a_315_75# 0.00121f
C89 VGND CIN 0.13789f
C90 VGND a_217_368# 0.0017f
C91 a_916_347# a_465_249# 0.0195f
C92 a_318_389# a_69_260# 0.02061f
C93 a_916_347# a_509_347# 0
C94 SUM B 0
C95 A a_69_260# 0.27191f
C96 a_465_249# a_1107_347# 0.15034f
C97 A VPB 0.14325f
C98 a_1107_347# COUT 0
C99 B CIN 0.19591f
C100 A a_237_75# 0.00252f
C101 a_936_75# A 0.00492f
C102 a_1100_75# a_69_260# 0
C103 VGND VNB 0.99802f
C104 COUT VNB 0.11284f
C105 CIN VNB 0.31573f
C106 A VNB 0.49885f
C107 VPWR VNB 0.79012f
C108 SUM VNB 0.11694f
C109 B VNB 0.61239f
C110 VPB VNB 2.08861f
C111 a_1100_75# VNB 0.01137f
C112 a_501_75# VNB 0.00504f
C113 a_1107_347# VNB 0.00204f
C114 a_509_347# VNB 0.00129f
C115 a_465_249# VNB 0.30402f
C116 a_69_260# VNB 0.15472f
.ends

.subckt sky130_fd_sc_hd__inv_8 a_60_47# w_n38_261# a_60_297# a_112_21# a_142_47# VSUBS
X0 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.16625 pd=1.5825 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16625 ps=1.5825 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10806 ps=1.145 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X3 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10806 ps=1.145 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X4 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.16625 pd=1.5825 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X5 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16625 ps=1.5825 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X6 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10806 ps=1.145 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X7 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.16625 pd=1.5825 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X8 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10806 ps=1.145 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X9 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16625 ps=1.5825 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X10 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.16625 pd=1.5825 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X11 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.10806 pd=1.145 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X12 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.10806 pd=1.145 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X13 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.10806 pd=1.145 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X14 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16625 ps=1.5825 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X15 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.10806 pd=1.145 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
C0 w_n38_261# a_60_47# 0.00793f
C1 a_60_47# a_142_47# 0.5745f
C2 w_n38_261# a_142_47# 0.03479f
C3 a_60_297# a_60_47# 0.08543f
C4 w_n38_261# a_60_297# 0.10021f
C5 a_60_47# a_112_21# 0.11686f
C6 a_60_297# a_142_47# 0.77995f
C7 w_n38_261# a_112_21# 0.25409f
C8 a_112_21# a_142_47# 0.82932f
C9 a_60_297# a_112_21# 0.12758f
C10 a_60_47# VSUBS 0.51049f
C11 a_142_47# VSUBS 0.12674f
C12 a_60_297# VSUBS 0.44991f
C13 a_112_21# VSUBS 0.77126f
C14 w_n38_261# VSUBS 0.87055f
.ends

.subckt sky130_fd_sc_hd__inv_12 a_60_47# w_n38_261# a_60_297# a_112_21# a_142_47#
+ VSUBS
X0 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.17708 pd=1.52083 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17708 ps=1.52083 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17708 ps=1.52083 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.17708 pd=1.52083 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=20600,606
X4 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1151 ps=1.1125 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X5 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1151 ps=1.1125 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.17708 pd=1.52083 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X7 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.17708 pd=1.52083 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1151 ps=1.1125 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X9 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1151 ps=1.1125 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X10 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17708 ps=1.52083 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X11 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1151 pd=1.1125 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=13390,466
X12 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1151 pd=1.1125 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X13 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17708 ps=1.52083 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X14 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1151 ps=1.1125 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X15 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.17708 pd=1.52083 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X16 a_142_47# a_112_21# a_60_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1151 ps=1.1125 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X17 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17708 ps=1.52083 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X18 a_60_297# a_112_21# a_142_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.17708 pd=1.52083 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X19 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1151 pd=1.1125 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X20 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1151 pd=1.1125 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X21 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1151 pd=1.1125 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X22 a_142_47# a_112_21# a_60_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17708 ps=1.52083 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X23 a_60_47# a_112_21# a_142_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1151 pd=1.1125 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 w_n38_261# a_60_47# 0.00933f
C1 a_60_47# a_142_47# 0.84337f
C2 w_n38_261# a_142_47# 0.04034f
C3 a_60_297# a_60_47# 0.12412f
C4 w_n38_261# a_60_297# 0.13063f
C5 a_60_47# a_112_21# 0.1674f
C6 a_60_297# a_142_47# 1.14598f
C7 w_n38_261# a_112_21# 0.38347f
C8 a_112_21# a_142_47# 1.26141f
C9 a_60_297# a_112_21# 0.18175f
C10 a_60_47# VSUBS 0.69459f
C11 a_142_47# VSUBS 0.13281f
C12 a_60_297# VSUBS 0.60586f
C13 a_112_21# VSUBS 1.13688f
C14 w_n38_261# VSUBS 1.22494f
.ends

.subckt sky130_fd_sc_hd__inv_6 a_37_47# w_n38_261# a_27_297# a_143_47# a_21_199# VSUBS
X0 a_27_297# a_21_199# a_143_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.20667 pd=1.74667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X1 a_143_47# a_21_199# a_27_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20667 ps=1.74667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 a_143_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12892 ps=1.26333 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X3 a_27_297# a_21_199# a_143_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.20667 pd=1.74667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 a_143_47# a_21_199# a_27_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20667 ps=1.74667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X5 a_27_297# a_21_199# a_143_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.20667 pd=1.74667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X6 a_143_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12892 ps=1.26333 w=0.65 l=0.15
**devattr s=9880,412 d=3510,184
X7 a_143_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12892 ps=1.26333 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X8 a_143_47# a_21_199# a_27_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20667 ps=1.74667 w=1 l=0.15
**devattr s=17200,572 d=5400,254
X9 a_37_47# a_21_199# a_143_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12892 pd=1.26333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X10 a_37_47# a_21_199# a_143_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12892 pd=1.26333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X11 a_37_47# a_21_199# a_143_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12892 pd=1.26333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=7020,368
C0 w_n38_261# a_37_47# 0.00676f
C1 a_37_47# a_143_47# 0.32587f
C2 w_n38_261# a_143_47# 0.01838f
C3 a_27_297# a_37_47# 0.06953f
C4 w_n38_261# a_27_297# 0.07832f
C5 a_37_47# a_21_199# 0.1215f
C6 a_27_297# a_143_47# 0.53032f
C7 w_n38_261# a_21_199# 0.21261f
C8 a_21_199# a_143_47# 0.54356f
C9 a_27_297# a_21_199# 0.13608f
C10 a_37_47# VSUBS 0.42142f
C11 a_143_47# VSUBS 0.09005f
C12 a_27_297# VSUBS 0.37325f
C13 a_21_199# VSUBS 0.64634f
C14 w_n38_261# VSUBS 0.69336f
.ends

.subckt sky130_fd_sc_hd__inv_4 a_37_47# w_n38_261# a_37_297# a_119_47# a_21_199# VSUBS
X0 a_37_297# a_21_199# a_119_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 a_119_47# a_21_199# a_37_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 a_119_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12837 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_37_297# a_21_199# a_119_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 a_37_47# a_21_199# a_119_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12837 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X5 a_119_47# a_21_199# a_37_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X6 a_37_47# a_21_199# a_119_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.12837 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X7 a_119_47# a_21_199# a_37_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12837 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 w_n38_261# a_37_47# 0.00667f
C1 a_37_47# a_119_47# 0.26259f
C2 w_n38_261# a_119_47# 0.0159f
C3 a_37_297# a_37_47# 0.05009f
C4 w_n38_261# a_37_297# 0.06539f
C5 a_37_47# a_21_199# 0.08191f
C6 a_37_297# a_119_47# 0.36178f
C7 w_n38_261# a_21_199# 0.14198f
C8 a_21_199# a_119_47# 0.35989f
C9 a_37_297# a_21_199# 0.09823f
C10 a_37_47# VSUBS 0.32682f
C11 a_119_47# VSUBS 0.08495f
C12 a_37_297# VSUBS 0.29639f
C13 a_21_199# VSUBS 0.45186f
C14 w_n38_261# VSUBS 0.51617f
.ends

.subckt sky130_fd_sc_hd__inv_2 w_n38_261# a_111_47# a_29_47# a_21_199# a_29_297# VSUBS
X0 a_111_47# a_21_199# a_29_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1 a_29_47# a_21_199# a_111_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 a_111_47# a_21_199# a_29_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_29_297# a_21_199# a_111_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
C0 w_n38_261# a_29_47# 0.00649f
C1 a_29_47# a_111_47# 0.1546f
C2 w_n38_261# a_111_47# 0.0061f
C3 a_29_297# a_29_47# 0.04227f
C4 w_n38_261# a_29_297# 0.05206f
C5 a_29_47# a_21_199# 0.06375f
C6 a_29_297# a_111_47# 0.2091f
C7 w_n38_261# a_21_199# 0.07418f
C8 a_21_199# a_111_47# 0.08939f
C9 a_29_297# a_21_199# 0.06305f
C10 a_29_47# VSUBS 0.26619f
C11 a_111_47# VSUBS 0.03316f
C12 a_29_297# VSUBS 0.24604f
C13 a_21_199# VSUBS 0.26281f
C14 w_n38_261# VSUBS 0.33898f
.ends

.subckt sky130_fd_sc_hs__inv_2 a_114_368# w_n38_332# a_27_368# a_30_74# a_21_260#
+ VSUBS
X0 a_114_368# a_21_260# a_30_74# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
**devattr s=8436,410 d=4144,204
X1 a_27_368# a_21_260# a_114_368# w_n38_332# sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
**devattr s=6720,284 d=12768,562
X2 a_30_74# a_21_260# a_114_368# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
**devattr s=4144,204 d=8436,410
X3 a_114_368# a_21_260# a_27_368# w_n38_332# sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
**devattr s=12768,562 d=6720,284
C0 w_n38_332# a_30_74# 0.00523f
C1 a_30_74# a_114_368# 0.16424f
C2 w_n38_332# a_114_368# 0.00641f
C3 a_27_368# a_30_74# 0.0376f
C4 w_n38_332# a_27_368# 0.06315f
C5 a_30_74# a_21_260# 0.06173f
C6 a_27_368# a_114_368# 0.21165f
C7 w_n38_332# a_21_260# 0.07759f
C8 a_21_260# a_114_368# 0.11388f
C9 a_27_368# a_21_260# 0.07533f
C10 a_30_74# VSUBS 0.30324f
C11 a_114_368# VSUBS 0.04146f
C12 a_27_368# VSUBS 0.26758f
C13 a_21_260# VSUBS 0.30548f
C14 w_n38_332# VSUBS 0.40622f
.ends

.subckt sky130_fd_sc_hd__inv_16 a_40_297# w_n38_261# a_40_47# a_26_199# a_122_47#
+ VSUBS
X0 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X2 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X3 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X5 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X7 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X8 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X10 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X11 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X12 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X13 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X14 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X15 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X16 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X17 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X18 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X19 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X20 a_40_47# a_26_199# a_122_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.09791 pd=1.0325 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X21 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X22 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X23 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X24 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X25 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X26 a_122_47# a_26_199# a_40_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15063 ps=1.42625 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X27 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X28 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X29 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X30 a_40_297# a_26_199# a_122_47# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.15063 pd=1.42625 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X31 a_122_47# a_26_199# a_40_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09791 ps=1.0325 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 w_n38_261# a_40_47# 0.01319f
C1 a_40_47# a_122_47# 1.06261f
C2 w_n38_261# a_122_47# 0.03049f
C3 a_40_297# a_40_47# 0.16076f
C4 w_n38_261# a_40_297# 0.15932f
C5 a_40_47# a_26_199# 0.26587f
C6 a_40_297# a_122_47# 1.46621f
C7 w_n38_261# a_26_199# 0.52574f
C8 a_26_199# a_122_47# 1.4347f
C9 a_40_297# a_26_199# 0.28026f
C10 a_40_47# VSUBS 0.86454f
C11 a_122_47# VSUBS 0.05506f
C12 a_40_297# VSUBS 0.73707f
C13 a_26_199# VSUBS 1.54575f
C14 w_n38_261# VSUBS 1.49072f
.ends

.subckt sky130_fd_sc_hd__inv_1 a_150_47# w_n38_261# a_68_47# a_68_297# a_64_199# VSUBS
X0 a_150_47# a_64_199# a_68_47# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1 a_150_47# a_64_199# a_68_297# w_n38_261# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
C0 w_n38_261# a_68_47# 0.00948f
C1 a_68_47# a_150_47# 0.09984f
C2 w_n38_261# a_150_47# 0.01774f
C3 a_68_297# a_68_47# 0.03382f
C4 w_n38_261# a_68_297# 0.05448f
C5 a_68_47# a_64_199# 0.04004f
C6 a_68_297# a_150_47# 0.12758f
C7 w_n38_261# a_64_199# 0.04506f
C8 a_64_199# a_150_47# 0.0476f
C9 a_68_297# a_64_199# 0.03703f
C10 a_68_47# VSUBS 0.25113f
C11 a_150_47# VSUBS 0.0961f
C12 a_68_297# VSUBS 0.21892f
C13 a_64_199# VSUBS 0.16664f
C14 w_n38_261# VSUBS 0.33898f
.ends

.subckt tt_um_ohmy90_ringOscillator clk A B CIN ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
Xsky130_fd_sc_hs__fa_1_6 A B sky130_fd_sc_hs__fa_1_6/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_4/CIN
+ SUM a_12918_2677# a_12925_2949# a_12136_2991# a_12133_2677# a_12734_2949# a_11902_3194#
+ a_12754_2677# a_13432_3194# a_12055_2677# a_12319_2677# a_12327_2949# a_12035_2970#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_7 A B sky130_fd_sc_hs__fa_1_7/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_6/CIN
+ SUM a_10856_2681# a_10863_2953# a_10074_2995# a_10071_2681# a_10672_2953# a_9840_3198#
+ a_10692_2681# a_11370_3198# a_9993_2681# a_10257_2681# a_10265_2953# a_9973_2974#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hd__inv_8_0 A sky130_fd_sc_hd__inv_8_0/w_n38_261# B li_21382_2780# li_22548_2776#
+ VNB sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__inv_12_0 A sky130_fd_sc_hd__inv_12_0/w_n38_261# B li_22548_2776#
+ li_24080_2768# VNB sky130_fd_sc_hd__inv_12
Xsky130_fd_sc_hd__inv_6_0 A sky130_fd_sc_hd__inv_6_0/w_n38_261# B li_21382_2780# COUT
+ VNB sky130_fd_sc_hd__inv_6
Xsky130_fd_sc_hd__inv_4_0 A sky130_fd_sc_hd__inv_4_0/w_n38_261# B COUT COUT VNB sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/w_n38_261# COUT A COUT B VNB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hs__fa_1_0 A B CIN A VNB VPB B sky130_fd_sc_hs__fa_1_1/CIN SUM a_2598_2695#
+ a_2605_2967# a_1816_3009# a_1813_2695# a_2414_2967# a_1582_3212# a_2434_2695# a_3112_3212#
+ a_1735_2695# a_1999_2695# a_2007_2967# a_1715_2988# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__inv_2_0 CIN sky130_fd_sc_hs__inv_2_0/w_n38_332# B A COUT VNB sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__fa_1_1 A B sky130_fd_sc_hs__fa_1_1/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_3/CIN
+ SUM a_4660_2691# a_4667_2963# a_3878_3005# a_3875_2691# a_4476_2963# a_3644_3208#
+ a_4496_2691# a_5174_3208# a_3797_2691# a_4061_2691# a_4069_2963# a_3777_2984# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hd__inv_16_0 B sky130_fd_sc_hd__inv_16_0/w_n38_261# A li_24080_2768#
+ a_27644_3049# VNB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_1_0 COUT sky130_fd_sc_hd__inv_1_0/w_n38_261# A B COUT VNB sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 COUT w_18084_2861# A B COUT VNB sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hs__fa_1_2 A B sky130_fd_sc_hs__fa_1_2/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_7/CIN
+ SUM a_8796_2685# a_8803_2957# a_8014_2999# a_8011_2685# a_8612_2957# a_7780_3202#
+ a_8632_2685# a_9310_3202# a_7933_2685# a_8197_2685# a_8205_2957# a_7913_2978# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hd__inv_16_1 B w_26254_2813# A a_27644_3049# a_29450_3031# VNB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hs__fa_1_4 A B sky130_fd_sc_hs__fa_1_4/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_5/CIN
+ SUM a_14992_2675# a_14999_2947# a_14210_2989# a_14207_2675# a_14808_2947# a_13976_3192#
+ a_14828_2675# a_15506_3192# a_14129_2675# a_14393_2675# a_14401_2947# a_14109_2968#
+ sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hs__fa_1_3 A B sky130_fd_sc_hs__fa_1_3/CIN A VNB VPB B sky130_fd_sc_hs__fa_1_2/CIN
+ SUM a_6734_2689# a_6741_2961# a_5952_3003# a_5949_2689# a_6550_2961# a_5718_3206#
+ a_6570_2689# a_7248_3206# a_5871_2689# a_6135_2689# a_6143_2961# a_5851_2982# sky130_fd_sc_hs__fa_1
Xsky130_fd_sc_hd__inv_16_2 B w_28060_2795# A a_29450_3031# ua[0] VNB sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hs__fa_1_5 A B sky130_fd_sc_hs__fa_1_5/CIN A VNB VPB B COUT SUM a_17054_2671#
+ a_17061_2943# a_16272_2985# a_16269_2671# a_16870_2943# a_16038_3188# a_16890_2671#
+ a_17568_3188# a_16191_2671# a_16455_2671# a_16463_2943# a_16171_2964# sky130_fd_sc_hs__fa_1
C0 a_3112_3212# a_1735_2695# 0
C1 a_14999_2947# sky130_fd_sc_hs__fa_1_5/CIN 0
C2 a_1999_2695# a_1582_3212# 0
C3 sky130_fd_sc_hs__fa_1_5/CIN a_16890_2671# -0
C4 uio_out[1] uio_out[0] 0.03102f
C5 a_10856_2681# a_9310_3202# 0
C6 B a_10074_2995# 0.00255f
C7 a_11902_3194# sky130_fd_sc_hs__fa_1_6/CIN 0.06636f
C8 a_5174_3208# a_4496_2691# -0
C9 B a_8014_2999# 0.00253f
C10 a_9310_3202# A 0.02705f
C11 sky130_fd_sc_hs__fa_1_7/CIN a_11370_3198# 0
C12 a_10265_2953# a_11370_3198# -0
C13 a_16191_2671# A 0
C14 a_12133_2677# A 0
C15 B a_8796_2685# 0.00714f
C16 a_8011_2685# A 0
C17 a_11902_3194# COUT 0.00172f
C18 a_10257_2681# a_11370_3198# 0
C19 sky130_fd_sc_hd__inv_6_0/w_n38_261# li_21382_2780# 0.00955f
C20 SUM a_7248_3206# 0
C21 a_2605_2967# sky130_fd_sc_hs__fa_1_1/CIN 0
C22 B a_8612_2957# 0.0053f
C23 sky130_fd_sc_hs__fa_1_6/CIN a_12918_2677# 0
C24 a_1813_2695# A 0.00102f
C25 sky130_fd_sc_hd__inv_8_0/w_n38_261# COUT 0
C26 li_22548_2776# a_27644_3049# 0
C27 B a_10863_2953# 0.05151f
C28 sky130_fd_sc_hs__fa_1_7/CIN a_9310_3202# 0.00636f
C29 B a_3112_3212# 0.0494f
C30 a_12918_2677# COUT 0
C31 B a_12055_2677# -0
C32 a_5851_2982# CIN 0
C33 a_9840_3198# COUT 0.00173f
C34 sky130_fd_sc_hs__fa_1_1/CIN a_4660_2691# 0
C35 VPB a_7248_3206# 0
C36 sky130_fd_sc_hs__fa_1_5/CIN sky130_fd_sc_hs__fa_1_4/CIN -0
C37 a_1816_3009# CIN 0.00257f
C38 a_6741_2961# sky130_fd_sc_hs__fa_1_3/CIN 0
C39 a_16038_3188# a_15506_3192# 0.00606f
C40 a_3112_3212# a_1582_3212# 0
C41 sky130_fd_sc_hs__fa_1_2/CIN a_7913_2978# 0.00449f
C42 a_13976_3192# a_15506_3192# -0
C43 a_14393_2675# sky130_fd_sc_hs__fa_1_4/CIN 0
C44 li_21382_2780# COUT 0.03717f
C45 sky130_fd_sc_hs__fa_1_5/CIN a_17061_2943# -0
C46 a_9310_3202# a_8205_2957# 0
C47 uo_out[3] uo_out[4] 0.03102f
C48 a_29450_3031# li_24080_2768# 0
C49 B a_4061_2691# 0.00186f
C50 B a_12319_2677# 0.00182f
C51 rst_n ui_in[0] 0.03102f
C52 a_10692_2681# B 0.00114f
C53 a_16272_2985# A 0
C54 A a_3777_2984# -0
C55 a_27644_3049# li_24080_2768# 0.04442f
C56 CIN a_3644_3208# 0.00209f
C57 CIN sky130_fd_sc_hs__fa_1_3/CIN 0.00252f
C58 B sky130_fd_sc_hd__inv_1_0/w_n38_261# 0.01732f
C59 B sky130_fd_sc_hs__fa_1_2/CIN 0.14387f
C60 a_16038_3188# A 0.00658f
C61 sky130_fd_sc_hs__fa_1_6/CIN a_11370_3198# 0.00642f
C62 B a_9993_2681# -0
C63 B a_12754_2677# 0.00113f
C64 a_11902_3194# SUM 0
C65 a_13976_3192# a_13432_3194# 0.00609f
C66 a_13976_3192# A 0.00662f
C67 a_12925_2949# B 0.05134f
C68 sky130_fd_sc_hs__fa_1_2/CIN a_7780_3202# 0.06636f
C69 a_5949_2689# CIN 0
C70 a_11370_3198# COUT 0.00229f
C71 sky130_fd_sc_hs__fa_1_5/CIN COUT 0.00486f
C72 a_11902_3194# VPB 0
C73 A a_6741_2961# 0
C74 uo_out[7] uio_out[0] 0.03102f
C75 a_17568_3188# sky130_fd_sc_hs__fa_1_5/CIN 0
C76 a_13976_3192# a_14207_2675# 0
C77 a_6734_2689# sky130_fd_sc_hs__fa_1_2/CIN -0
C78 a_14393_2675# COUT 0
C79 SUM a_9840_3198# 0
C80 B a_16455_2671# 0.0018f
C81 a_6570_2689# sky130_fd_sc_hs__fa_1_3/CIN -0
C82 a_5851_2982# sky130_fd_sc_hs__fa_1_3/CIN 0.0045f
C83 CIN a_3797_2691# 0
C84 B a_2605_2967# 0.05291f
C85 li_22548_2776# sky130_fd_sc_hd__inv_16_0/w_n38_261# 0.0011f
C86 a_12133_2677# sky130_fd_sc_hs__fa_1_6/CIN 0
C87 a_3112_3212# a_2598_2695# -0
C88 CIN A 0.21476f
C89 a_2434_2695# a_3112_3212# 0
C90 a_9310_3202# COUT 0.00204f
C91 a_16191_2671# COUT 0
C92 VPB a_9840_3198# 0
C93 li_24080_2768# w_26254_2813# 0
C94 a_12133_2677# COUT 0
C95 B a_4660_2691# 0.00758f
C96 a_16171_2964# A -0
C97 B a_14210_2989# 0.00249f
C98 B a_2414_2967# 0.00514f
C99 B a_7248_3206# 0.04438f
C100 A sky130_fd_sc_hd__inv_2_0/w_n38_261# 0
C101 a_4496_2691# sky130_fd_sc_hs__fa_1_1/CIN -0
C102 A a_14129_2675# 0
C103 a_2007_2967# a_3112_3212# -0
C104 B a_7933_2685# -0
C105 sky130_fd_sc_hd__inv_16_0/w_n38_261# li_24080_2768# 0.00978f
C106 a_13976_3192# sky130_fd_sc_hs__fa_1_4/CIN 0.06234f
C107 a_7780_3202# a_7248_3206# 0.00606f
C108 a_13976_3192# a_14109_2968# -0
C109 a_5949_2689# sky130_fd_sc_hs__fa_1_3/CIN 0
C110 a_3112_3212# a_1999_2695# -0
C111 SUM a_11370_3198# 0
C112 a_6570_2689# A 0.0048f
C113 B a_16463_2943# 0.00626f
C114 li_22548_2776# B 0.13535f
C115 a_5851_2982# A -0
C116 a_5718_3206# a_7248_3206# 0
C117 sky130_fd_sc_hs__fa_1_5/CIN SUM 0.07889f
C118 B sky130_fd_sc_hs__inv_2_0/w_n38_332# 0.01636f
C119 a_1816_3009# A 0.00186f
C120 sky130_fd_sc_hs__fa_1_2/CIN a_8197_2685# 0
C121 clk rst_n 0.03102f
C122 a_16269_2671# A 0
C123 CIN a_5871_2689# 0
C124 a_6734_2689# a_7248_3206# -0
C125 CIN a_8205_2957# 0
C126 VPB a_11370_3198# 0.00733f
C127 a_9973_2974# A -0
C128 li_21382_2780# sky130_fd_sc_hd__inv_4_0/w_n38_261# 0
C129 B a_5952_3003# 0.00251f
C130 VPB sky130_fd_sc_hs__fa_1_5/CIN 0.02471f
C131 A a_3644_3208# 0.05984f
C132 A sky130_fd_sc_hs__fa_1_3/CIN 0.14599f
C133 a_16272_2985# COUT 0
C134 a_9310_3202# SUM 0
C135 B a_14828_2675# 0.00115f
C136 A a_12734_2949# 0.0028f
C137 a_12734_2949# a_13432_3194# 0
C138 a_5174_3208# CIN 0.0025f
C139 a_11902_3194# B 0.00724f
C140 li_22548_2776# sky130_fd_sc_hd__inv_12_0/w_n38_261# 0.00918f
C141 a_16038_3188# COUT 0.00208f
C142 ui_in[7] uio_in[0] 0.03102f
C143 B li_24080_2768# 0.13983f
C144 a_17568_3188# a_16038_3188# 0
C145 a_13976_3192# COUT 0.00174f
C146 sky130_fd_sc_hs__fa_1_2/CIN a_8014_2999# 0
C147 CIN a_6143_2961# 0
C148 a_5949_2689# A 0
C149 B sky130_fd_sc_hd__inv_8_0/w_n38_261# 0.01204f
C150 VPB a_9310_3202# 0
C151 a_9973_2974# sky130_fd_sc_hs__fa_1_7/CIN 0.00447f
C152 sky130_fd_sc_hs__fa_1_4/CIN a_14129_2675# 0.00124f
C153 a_15506_3192# A 0.0316f
C154 a_8796_2685# sky130_fd_sc_hs__fa_1_2/CIN 0
C155 CIN a_3875_2691# 0
C156 B a_12918_2677# 0.0071f
C157 B a_9840_3198# 0.00738f
C158 B a_4496_2691# 0.00114f
C159 sky130_fd_sc_hs__fa_1_2/CIN a_8612_2957# 0
C160 sky130_fd_sc_hd__inv_12_0/w_n38_261# li_24080_2768# 0.00547f
C161 a_3797_2691# A 0.00203f
C162 a_6550_2961# sky130_fd_sc_hs__fa_1_3/CIN 0
C163 B li_21382_2780# 0.14494f
C164 a_10856_2681# A 0.01142f
C165 CIN a_4069_2963# 0.00118f
C166 A a_13432_3194# 0.03092f
C167 a_5871_2689# sky130_fd_sc_hs__fa_1_3/CIN 0.00124f
C168 a_10071_2681# a_9840_3198# 0
C169 CIN COUT 0.09476f
C170 a_16171_2964# COUT 0
C171 B a_6135_2689# 0.00209f
C172 a_14999_2947# A 0
C173 a_16890_2671# A 0.00477f
C174 a_5174_3208# a_3644_3208# 0
C175 a_5174_3208# sky130_fd_sc_hs__fa_1_3/CIN 0.00595f
C176 a_16038_3188# SUM 0
C177 COUT sky130_fd_sc_hd__inv_2_0/w_n38_261# 0.019f
C178 a_14129_2675# COUT 0
C179 A a_14207_2675# 0
C180 li_21382_2780# sky130_fd_sc_hd__inv_12_0/w_n38_261# 0.00111f
C181 a_12035_2970# A -0
C182 a_10856_2681# sky130_fd_sc_hs__fa_1_7/CIN 0
C183 a_13976_3192# SUM 0
C184 B a_11370_3198# 0.04956f
C185 uo_out[0] uio_in[7] 0.03102f
C186 sky130_fd_sc_hs__fa_1_7/CIN A 0.14708f
C187 a_6143_2961# sky130_fd_sc_hs__fa_1_3/CIN 0
C188 a_8632_2685# A 0.00477f
C189 a_10265_2953# A 0.00223f
C190 a_5718_3206# a_6135_2689# 0
C191 B sky130_fd_sc_hs__fa_1_5/CIN 0.12687f
C192 A w_28060_2795# 0.00308f
C193 a_3777_2984# sky130_fd_sc_hs__fa_1_1/CIN 0.00449f
C194 a_4476_2963# A 0.00282f
C195 a_16870_2943# sky130_fd_sc_hs__fa_1_5/CIN 0
C196 a_16038_3188# VPB 0
C197 a_15506_3192# sky130_fd_sc_hs__fa_1_4/CIN 0
C198 a_8796_2685# a_7248_3206# 0
C199 a_6550_2961# A 0.00288f
C200 B a_14393_2675# 0.00181f
C201 sky130_fd_sc_hs__fa_1_5/CIN a_17054_2671# 0
C202 a_10257_2681# A 0.00859f
C203 a_13976_3192# VPB 0
C204 A a_5871_2689# 0
C205 a_16269_2671# COUT 0
C206 A a_8205_2957# 0.00293f
C207 sky130_fd_sc_hs__fa_1_6/CIN a_12734_2949# 0
C208 a_9973_2974# COUT 0
C209 uio_in[3] uio_in[2] 0.03102f
C210 a_17568_3188# a_16269_2671# 0
C211 B a_9310_3202# 0.04713f
C212 a_3112_3212# a_4660_2691# 0
C213 sky130_fd_sc_hs__fa_1_7/CIN a_10265_2953# 0
C214 B a_16191_2671# -0
C215 CIN SUM 0.0047f
C216 B a_12133_2677# 0
C217 sky130_fd_sc_hs__fa_1_4/CIN a_13432_3194# 0.00595f
C218 sky130_fd_sc_hs__fa_1_4/CIN A 0.14323f
C219 a_5174_3208# A 0.03356f
C220 a_4667_2963# CIN 0
C221 A a_14109_2968# -0
C222 B a_8011_2685# 0
C223 a_9310_3202# a_7780_3202# 0
C224 A a_8803_2957# 0
C225 a_10257_2681# sky130_fd_sc_hs__fa_1_7/CIN 0
C226 A a_17061_2943# 0
C227 A a_6143_2961# 0.00252f
C228 A a_12327_2949# 0.00224f
C229 a_13432_3194# a_12327_2949# 0
C230 sky130_fd_sc_hd__inv_6_0/w_n38_261# A 0.00176f
C231 a_14999_2947# sky130_fd_sc_hs__fa_1_4/CIN 0
C232 B a_1813_2695# 0
C233 VPB CIN 0.0286f
C234 CIN sky130_fd_sc_hs__fa_1_1/CIN 0.00358f
C235 sky130_fd_sc_hs__fa_1_4/CIN a_14207_2675# 0
C236 a_15506_3192# COUT 0.00247f
C237 a_1813_2695# a_1582_3212# 0
C238 a_3875_2691# A 0.00209f
C239 a_10856_2681# sky130_fd_sc_hs__fa_1_6/CIN -0
C240 sky130_fd_sc_hs__fa_1_2/CIN a_7248_3206# 0.00578f
C241 sky130_fd_sc_hs__fa_1_6/CIN a_13432_3194# 0
C242 sky130_fd_sc_hs__fa_1_6/CIN A 0.14275f
C243 sky130_fd_sc_hs__fa_1_2/CIN a_7933_2685# 0.00126f
C244 a_5174_3208# a_4476_2963# -0
C245 sky130_fd_sc_hs__fa_1_7/CIN a_8803_2957# 0
C246 a_10856_2681# COUT 0
C247 a_4069_2963# A 0.0022f
C248 a_13432_3194# COUT 0.00233f
C249 A COUT 0.73879f
C250 ui_in[7] ui_in[6] 0.03102f
C251 ua[0] A 0.11504f
C252 B a_3777_2984# 0.00247f
C253 B a_16272_2985# 0.00251f
C254 a_17568_3188# A 0.0311f
C255 a_12035_2970# sky130_fd_sc_hs__fa_1_6/CIN 0.00449f
C256 SUM a_3644_3208# 0
C257 SUM sky130_fd_sc_hs__fa_1_3/CIN 0.07548f
C258 B a_16038_3188# 0.00717f
C259 uio_oe[0] uio_oe[1] 0.03102f
C260 a_14999_2947# COUT 0
C261 sky130_fd_sc_hs__fa_1_7/CIN sky130_fd_sc_hs__fa_1_6/CIN -0
C262 a_16890_2671# COUT 0
C263 a_4667_2963# sky130_fd_sc_hs__fa_1_3/CIN 0
C264 uio_out[1] uio_out[2] 0.03102f
C265 sky130_fd_sc_hs__fa_1_4/CIN a_14109_2968# 0.0045f
C266 B a_13976_3192# 0.00726f
C267 a_14207_2675# COUT 0
C268 CIN a_1715_2988# 0.0017f
C269 a_17568_3188# a_16890_2671# -0
C270 a_12035_2970# COUT 0
C271 sky130_fd_sc_hs__fa_1_7/CIN COUT 0.00278f
C272 VPB a_3644_3208# 0
C273 a_10265_2953# COUT 0.00105f
C274 VPB sky130_fd_sc_hs__fa_1_3/CIN 0.01875f
C275 a_15506_3192# SUM 0
C276 a_3644_3208# sky130_fd_sc_hs__fa_1_1/CIN 0.06636f
C277 sky130_fd_sc_hs__fa_1_1/CIN sky130_fd_sc_hs__fa_1_3/CIN -0
C278 B a_6741_2961# 0.05141f
C279 a_9310_3202# a_8197_2685# 0
C280 a_29450_3031# A 0.19868f
C281 ua[0] w_28060_2795# 0.00869f
C282 CIN a_7913_2978# 0
C283 a_27644_3049# A 0.19465f
C284 a_10257_2681# COUT 0
C285 sky130_fd_sc_hs__fa_1_6/CIN sky130_fd_sc_hs__fa_1_4/CIN -0
C286 COUT a_8205_2957# 0
C287 a_15506_3192# VPB 0
C288 B CIN 0.62951f
C289 SUM a_13432_3194# 0
C290 SUM A 0.02098f
C291 a_5174_3208# a_4069_2963# 0
C292 a_4667_2963# A 0
C293 sky130_fd_sc_hs__fa_1_6/CIN a_12327_2949# 0
C294 sky130_fd_sc_hs__fa_1_4/CIN COUT 0.00281f
C295 B a_16171_2964# 0.00245f
C296 CIN a_1582_3212# 0.00855f
C297 a_14109_2968# COUT 0
C298 CIN a_7780_3202# 0.00188f
C299 ui_in[4] ui_in[5] 0.03102f
C300 B sky130_fd_sc_hd__inv_2_0/w_n38_261# 0.01139f
C301 B a_14129_2675# -0
C302 a_29450_3031# w_28060_2795# 0.01123f
C303 a_8803_2957# COUT 0
C304 a_17061_2943# COUT 0.00339f
C305 a_5718_3206# CIN 0.00192f
C306 uio_in[3] uio_in[4] 0.03102f
C307 a_3797_2691# sky130_fd_sc_hs__fa_1_1/CIN 0.00126f
C308 a_12327_2949# COUT 0.00105f
C309 a_8796_2685# a_9310_3202# -0
C310 VPB a_13432_3194# 0
C311 VPB A 0.0505f
C312 a_27644_3049# w_28060_2795# 0.00158f
C313 sky130_fd_sc_hd__inv_6_0/w_n38_261# COUT 0.01373f
C314 A sky130_fd_sc_hs__fa_1_1/CIN 0.14974f
C315 a_6734_2689# CIN 0
C316 sky130_fd_sc_hs__fa_1_7/CIN SUM 0.07963f
C317 B a_6570_2689# 0.00111f
C318 a_9310_3202# a_8612_2957# -0
C319 B a_5851_2982# 0.00243f
C320 A w_18084_2861# 0.00133f
C321 a_1816_3009# B 0.00201f
C322 sky130_fd_sc_hs__fa_1_6/CIN COUT 0.0029f
C323 A w_26254_2813# 0.00298f
C324 B a_16269_2671# 0
C325 a_14808_2947# A 0.00282f
C326 uio_out[4] uio_out[5] 0.03102f
C327 B a_9973_2974# 0.00246f
C328 VPB sky130_fd_sc_hs__fa_1_7/CIN 0.01776f
C329 A sky130_fd_sc_hd__inv_4_0/w_n38_261# -0.00174f
C330 a_3878_3005# CIN 0
C331 a_10672_2953# A 0.00282f
C332 B a_3644_3208# 0.0075f
C333 B sky130_fd_sc_hs__fa_1_3/CIN 0.15242f
C334 a_17568_3188# COUT 0.02908f
C335 sky130_fd_sc_hd__inv_16_0/w_n38_261# A 0.00277f
C336 A a_1735_2695# 0
C337 B a_12734_2949# 0.00529f
C338 a_4476_2963# sky130_fd_sc_hs__fa_1_1/CIN 0
C339 li_22548_2776# li_24080_2768# 0.11802f
C340 SUM sky130_fd_sc_hs__fa_1_4/CIN 0.07548f
C341 a_5174_3208# SUM 0
C342 CIN a_2598_2695# 0
C343 uio_oe[5] uio_oe[6] 0.03102f
C344 a_1813_2695# a_3112_3212# -0
C345 a_2434_2695# CIN -0
C346 li_22548_2776# sky130_fd_sc_hd__inv_8_0/w_n38_261# 0.00649f
C347 A a_1715_2988# 0.00175f
C348 a_9310_3202# sky130_fd_sc_hs__fa_1_2/CIN 0
C349 a_5949_2689# B 0
C350 a_5718_3206# sky130_fd_sc_hs__fa_1_3/CIN 0.06234f
C351 B a_15506_3192# 0.04767f
C352 VPB sky130_fd_sc_hs__fa_1_4/CIN 0.01878f
C353 a_5174_3208# VPB 0
C354 sky130_fd_sc_hs__fa_1_2/CIN a_8011_2685# 0
C355 sky130_fd_sc_hs__fa_1_7/CIN a_10672_2953# 0
C356 sky130_fd_sc_hs__fa_1_5/CIN a_16455_2671# 0
C357 CIN a_8197_2685# 0
C358 a_6734_2689# sky130_fd_sc_hs__fa_1_3/CIN 0
C359 uio_oe[2] uio_oe[1] 0.03102f
C360 a_5174_3208# sky130_fd_sc_hs__fa_1_1/CIN 0
C361 A a_7913_2978# -0
C362 a_15506_3192# a_17054_2671# 0
C363 ua[0] a_29450_3031# 0.03424f
C364 a_6135_2689# a_7248_3206# 0
C365 a_2007_2967# CIN 0.01499f
C366 li_22548_2776# li_21382_2780# 0.16918f
C367 ua[0] a_27644_3049# 0
C368 a_5718_3206# a_5949_2689# 0
C369 B a_3797_2691# -0
C370 A a_12136_2991# 0
C371 sky130_fd_sc_hs__fa_1_6/CIN SUM 0.07889f
C372 B a_10856_2681# 0.00722f
C373 uio_in[1] uio_in[0] 0.03102f
C374 CIN a_1999_2695# 0.00138f
C375 B a_13432_3194# 0.04883f
C376 B A 16.71954f
C377 sky130_fd_sc_hd__inv_8_0/w_n38_261# li_24080_2768# 0.00106f
C378 a_14808_2947# sky130_fd_sc_hs__fa_1_4/CIN 0
C379 a_16870_2943# A 0.00282f
C380 uio_in[6] uio_in[7] 0.03102f
C381 SUM COUT 0.00322f
C382 a_17054_2671# A 0.01045f
C383 a_1582_3212# A 0.01636f
C384 a_3875_2691# sky130_fd_sc_hs__fa_1_1/CIN 0
C385 A a_7780_3202# 0.00653f
C386 VPB sky130_fd_sc_hs__fa_1_6/CIN 0.01755f
C387 CIN a_8014_2999# 0
C388 uio_oe[3] uio_oe[4] 0.03102f
C389 ui_in[3] ui_in[2] 0.03102f
C390 B a_14999_2947# 0.05133f
C391 B a_16890_2671# 0.00113f
C392 a_10071_2681# A 0
C393 B a_14207_2675# 0
C394 a_5718_3206# A 0.00671f
C395 B a_12035_2970# 0.00246f
C396 li_21382_2780# li_24080_2768# 0
C397 VPB COUT 0.03925f
C398 a_4069_2963# sky130_fd_sc_hs__fa_1_1/CIN 0
C399 a_15506_3192# a_14992_2675# -0
C400 a_27644_3049# a_29450_3031# 0.0354f
C401 sky130_fd_sc_hd__inv_12_0/w_n38_261# A 0.00306f
C402 B sky130_fd_sc_hs__fa_1_7/CIN 0.12798f
C403 B a_8632_2685# 0.00114f
C404 sky130_fd_sc_hs__fa_1_5/CIN a_16463_2943# 0
C405 a_6734_2689# A 0.01194f
C406 B a_10265_2953# 0.00622f
C407 a_17568_3188# VPB -0
C408 li_21382_2780# sky130_fd_sc_hd__inv_8_0/w_n38_261# 0.01474f
C409 B w_28060_2795# 0.01299f
C410 B a_4476_2963# 0.00531f
C411 uio_in[1] uio_in[2] 0.03102f
C412 B a_6550_2961# 0.00524f
C413 w_18084_2861# COUT 0.03098f
C414 a_10257_2681# B 0.00183f
C415 uo_out[1] uo_out[0] 0.03102f
C416 a_10071_2681# sky130_fd_sc_hs__fa_1_7/CIN 0
C417 B a_5871_2689# -0
C418 ua[0] w_26254_2813# 0
C419 a_17568_3188# w_18084_2861# 0.00123f
C420 a_3112_3212# CIN 0.03133f
C421 a_14992_2675# a_13432_3194# 0
C422 a_11902_3194# a_11370_3198# 0.00606f
C423 a_14992_2675# A 0.01055f
C424 B a_8205_2957# 0.00624f
C425 a_15506_3192# a_14401_2947# -0
C426 a_3878_3005# A 0
C427 sky130_fd_sc_hs__fa_1_2/CIN a_6741_2961# 0
C428 sky130_fd_sc_hd__inv_4_0/w_n38_261# COUT 0.02089f
C429 B sky130_fd_sc_hs__fa_1_4/CIN 0.1342f
C430 B a_5174_3208# 0.04984f
C431 B a_14109_2968# 0.00241f
C432 uo_out[7] uo_out[6] 0.03102f
C433 uio_out[2] uio_out[3] 0.03102f
C434 CIN a_4061_2691# 0
C435 a_5718_3206# a_5871_2689# -0
C436 a_2598_2695# A 0.01263f
C437 B a_8803_2957# 0.05139f
C438 B a_17061_2943# 0.05166f
C439 a_2434_2695# A 0.005f
C440 a_12918_2677# a_11370_3198# 0
C441 B a_6143_2961# 0.00745f
C442 CIN sky130_fd_sc_hs__fa_1_2/CIN 0.00209f
C443 B a_12327_2949# 0.00619f
C444 A a_14401_2947# 0.00225f
C445 a_11370_3198# a_9840_3198# -0
C446 sky130_fd_sc_hd__inv_6_0/w_n38_261# B 0.01259f
C447 a_29450_3031# w_26254_2813# 0.00766f
C448 a_5718_3206# a_5174_3208# 0.00609f
C449 VPB SUM 0.01931f
C450 a_27644_3049# w_26254_2813# 0.00966f
C451 a_8197_2685# A 0.00902f
C452 B a_3875_2691# 0
C453 SUM sky130_fd_sc_hs__fa_1_1/CIN 0.07889f
C454 sky130_fd_sc_hs__fa_1_6/CIN a_12136_2991# 0
C455 a_4667_2963# sky130_fd_sc_hs__fa_1_1/CIN -0
C456 a_5174_3208# a_6734_2689# 0
C457 B sky130_fd_sc_hs__fa_1_6/CIN 0.12612f
C458 a_2007_2967# A 0.0037f
C459 a_13976_3192# a_14210_2989# -0
C460 sky130_fd_sc_hd__inv_16_0/w_n38_261# a_29450_3031# 0
C461 a_12136_2991# COUT 0
C462 a_1999_2695# A 0.00974f
C463 B a_4069_2963# 0.00628f
C464 a_9310_3202# a_9840_3198# 0.00608f
C465 a_27644_3049# sky130_fd_sc_hd__inv_16_0/w_n38_261# 0.00832f
C466 VPB sky130_fd_sc_hs__fa_1_1/CIN 0.01757f
C467 a_3112_3212# a_3644_3208# 0.00606f
C468 B COUT 1.22264f
C469 ua[0] B 0.07667f
C470 uio_out[6] uio_out[5] 0.03102f
C471 a_16870_2943# COUT 0
C472 sky130_fd_sc_hs__fa_1_4/CIN a_14992_2675# 0
C473 a_2605_2967# CIN 0.00353f
C474 B a_17568_3188# 0.04871f
C475 A a_10074_2995# 0
C476 a_17054_2671# COUT 0.00228f
C477 a_17568_3188# a_16870_2943# 0
C478 A a_8014_2999# 0
C479 uo_out[6] uo_out[5] 0.03102f
C480 a_10071_2681# COUT 0
C481 a_8796_2685# A 0.01048f
C482 CIN a_4660_2691# 0
C483 a_2414_2967# CIN 0.0025f
C484 sky130_fd_sc_hs__fa_1_2/CIN sky130_fd_sc_hs__fa_1_3/CIN -0
C485 sky130_fd_sc_hd__inv_12_0/w_n38_261# COUT 0
C486 CIN a_7248_3206# 0.0032f
C487 sky130_fd_sc_hs__fa_1_4/CIN a_14401_2947# 0
C488 A a_8612_2957# 0.00282f
C489 B a_29450_3031# 0.16679f
C490 CIN a_7933_2685# 0
C491 sky130_fd_sc_hs__fa_1_7/CIN a_10074_2995# 0
C492 a_10863_2953# A 0.00117f
C493 B a_27644_3049# 0.16844f
C494 a_3112_3212# A 0.03499f
C495 uio_oe[5] uio_oe[4] 0.03102f
C496 a_8796_2685# sky130_fd_sc_hs__fa_1_7/CIN -0
C497 A a_12055_2677# 0
C498 a_14992_2675# COUT 0
C499 a_16191_2671# sky130_fd_sc_hs__fa_1_5/CIN 0.00126f
C500 CIN sky130_fd_sc_hs__inv_2_0/w_n38_332# 0.00808f
C501 B SUM 0.02967f
C502 a_4667_2963# B 0.05256f
C503 a_12319_2677# a_13432_3194# 0
C504 a_12319_2677# A 0.0086f
C505 A a_4061_2691# 0.07073f
C506 a_6570_2689# a_7248_3206# 0
C507 a_5952_3003# CIN 0
C508 sky130_fd_sc_hs__fa_1_7/CIN a_10863_2953# -0
C509 SUM a_1582_3212# 0
C510 SUM a_7780_3202# 0
C511 a_10692_2681# A 0.00477f
C512 a_27644_3049# sky130_fd_sc_hd__inv_12_0/w_n38_261# 0
C513 sky130_fd_sc_hd__inv_1_0/w_n38_261# A 0.00126f
C514 sky130_fd_sc_hs__fa_1_2/CIN A 0.1457f
C515 a_14401_2947# COUT 0.00104f
C516 B VPB 0.39646f
C517 a_5718_3206# SUM 0
C518 A a_9993_2681# 0
C519 B sky130_fd_sc_hs__fa_1_1/CIN 0.14445f
C520 sky130_fd_sc_hs__fa_1_3/CIN a_4660_2691# 0
C521 A a_12754_2677# 0.00476f
C522 uio_out[4] uio_out[3] 0.03102f
C523 a_12925_2949# A 0
C524 VPB a_1582_3212# 0
C525 VPB a_7780_3202# 0
C526 a_8197_2685# COUT 0
C527 a_7248_3206# sky130_fd_sc_hs__fa_1_3/CIN 0
C528 B w_18084_2861# 0.01776f
C529 a_5718_3206# VPB 0
C530 B w_26254_2813# 0.01675f
C531 a_10692_2681# sky130_fd_sc_hs__fa_1_7/CIN -0
C532 B a_14808_2947# 0.00529f
C533 sky130_fd_sc_hs__fa_1_7/CIN sky130_fd_sc_hs__fa_1_2/CIN -0
C534 sky130_fd_sc_hs__fa_1_2/CIN a_8632_2685# -0
C535 a_16272_2985# sky130_fd_sc_hs__fa_1_5/CIN 0
C536 uio_in[5] uio_in[4] 0.03102f
C537 uio_in[6] uio_in[5] 0.03102f
C538 A a_16455_2671# 0.00863f
C539 sky130_fd_sc_hs__fa_1_7/CIN a_9993_2681# 0.00127f
C540 a_16038_3188# sky130_fd_sc_hs__fa_1_5/CIN 0.06636f
C541 B sky130_fd_sc_hd__inv_4_0/w_n38_261# 0.01192f
C542 a_2605_2967# A 0.00106f
C543 B a_10672_2953# 0.00529f
C544 ui_in[0] ui_in[1] 0.03102f
C545 B sky130_fd_sc_hd__inv_16_0/w_n38_261# 0.01669f
C546 B a_1735_2695# 0
C547 a_10074_2995# COUT 0
C548 a_13976_3192# a_14393_2675# 0
C549 sky130_fd_sc_hs__fa_1_2/CIN a_8205_2957# 0
C550 a_1582_3212# a_1735_2695# -0
C551 B a_1715_2988# 0.00185f
C552 A a_4660_2691# 0.01189f
C553 a_5952_3003# sky130_fd_sc_hs__fa_1_3/CIN 0
C554 a_8796_2685# COUT 0
C555 a_14210_2989# A 0
C556 CIN a_6135_2689# 0
C557 a_5174_3208# a_4061_2691# 0
C558 uio_oe[0] uio_out[7] 0.03102f
C559 a_2414_2967# A 0.00335f
C560 sky130_fd_sc_hs__fa_1_6/CIN a_10863_2953# 0
C561 A a_7248_3206# 0.02842f
C562 a_3878_3005# sky130_fd_sc_hs__fa_1_1/CIN 0
C563 ui_in[2] ui_in[1] 0.03102f
C564 A a_7933_2685# 0
C565 sky130_fd_sc_hs__fa_1_6/CIN a_12055_2677# 0.00126f
C566 B a_7913_2978# 0.00247f
C567 sky130_fd_sc_hs__fa_1_2/CIN a_8803_2957# -0
C568 a_12925_2949# sky130_fd_sc_hs__fa_1_4/CIN 0
C569 a_10863_2953# COUT 0
C570 ui_in[3] ui_in[4] 0.03102f
C571 uo_out[2] uo_out[3] 0.03102f
C572 a_2598_2695# sky130_fd_sc_hs__fa_1_1/CIN -0
C573 a_9973_2974# a_9840_3198# 0
C574 B a_12136_2991# 0.00252f
C575 li_22548_2776# A 0.15339f
C576 a_16463_2943# A 0.00226f
C577 a_12055_2677# COUT 0
C578 A sky130_fd_sc_hs__inv_2_0/w_n38_332# 0
C579 sky130_fd_sc_hs__fa_1_6/CIN a_12319_2677# 0
C580 uio_oe[3] uio_oe[2] 0.03102f
C581 sky130_fd_sc_hs__fa_1_5/CIN a_16171_2964# 0.00449f
C582 B a_16870_2943# 0.00543f
C583 B a_1582_3212# 0.01109f
C584 B a_17054_2671# 0.00708f
C585 B a_7780_3202# 0.00739f
C586 a_5952_3003# A 0
C587 a_12319_2677# COUT 0
C588 a_9310_3202# CIN 0
C589 B a_10071_2681# 0
C590 sky130_fd_sc_hs__fa_1_6/CIN a_12754_2677# -0
C591 uio_out[6] uio_out[7] 0.03102f
C592 a_12925_2949# sky130_fd_sc_hs__fa_1_6/CIN -0
C593 a_5718_3206# B 0.00747f
C594 a_14828_2675# A 0.00477f
C595 sky130_fd_sc_hd__inv_1_0/w_n38_261# COUT 0.02878f
C596 a_11902_3194# A 0.00651f
C597 a_11902_3194# a_13432_3194# 0
C598 sky130_fd_sc_hs__fa_1_2/CIN COUT 0
C599 CIN a_8011_2685# 0
C600 a_17568_3188# sky130_fd_sc_hd__inv_1_0/w_n38_261# 0
C601 B sky130_fd_sc_hd__inv_12_0/w_n38_261# 0.0156f
C602 uo_out[5] uo_out[4] 0.03102f
C603 a_9993_2681# COUT 0
C604 li_24080_2768# A 0.16193f
C605 a_6135_2689# sky130_fd_sc_hs__fa_1_3/CIN 0
C606 B a_6734_2689# 0.00716f
C607 a_5174_3208# a_4660_2691# -0
C608 a_14210_2989# sky130_fd_sc_hs__fa_1_4/CIN 0
C609 a_12925_2949# COUT 0
C610 sky130_fd_sc_hd__inv_8_0/w_n38_261# A 0.00107f
C611 a_16269_2671# sky130_fd_sc_hs__fa_1_5/CIN 0
C612 clk ena 0.03102f
C613 a_12918_2677# a_13432_3194# -0
C614 a_12918_2677# A 0.0105f
C615 uo_out[2] uo_out[1] 0.03102f
C616 A a_9840_3198# 0.00641f
C617 B a_14992_2675# 0.00709f
C618 a_7248_3206# a_6143_2961# -0
C619 a_3112_3212# SUM 0
C620 A a_4496_2691# 0.00523f
C621 a_16455_2671# COUT 0
C622 B a_3878_3005# 0.00253f
C623 li_21382_2780# A 0.15105f
C624 a_17568_3188# a_16455_2671# 0
C625 uio_oe[7] uio_oe[6] 0.03102f
C626 B a_2598_2695# 0.00768f
C627 ui_in[6] ui_in[5] 0.03102f
C628 VPB a_3112_3212# 0
C629 CIN a_3777_2984# 0
C630 sky130_fd_sc_hd__inv_6_0/w_n38_261# li_22548_2776# 0.00103f
C631 B a_2434_2695# 0.00116f
C632 a_15506_3192# sky130_fd_sc_hs__fa_1_5/CIN 0.00578f
C633 B a_14401_2947# 0.00607f
C634 a_3112_3212# sky130_fd_sc_hs__fa_1_1/CIN 0.00578f
C635 A a_6135_2689# 0.00862f
C636 a_14210_2989# COUT 0
C637 sky130_fd_sc_hs__fa_1_7/CIN a_9840_3198# 0.06628f
C638 sky130_fd_sc_hs__fa_1_2/CIN SUM 0.07889f
C639 a_15506_3192# a_14393_2675# 0
C640 a_14828_2675# sky130_fd_sc_hs__fa_1_4/CIN -0
C641 a_2434_2695# a_1582_3212# -0
C642 a_10856_2681# a_11370_3198# -0
C643 B a_8197_2685# 0.00184f
C644 A a_11370_3198# 0.03199f
C645 a_10257_2681# a_9840_3198# 0
C646 B a_2007_2967# 0.00539f
C647 a_4061_2691# sky130_fd_sc_hs__fa_1_1/CIN 0
C648 sky130_fd_sc_hs__fa_1_5/CIN A 0.14329f
C649 VPB sky130_fd_sc_hs__fa_1_2/CIN 0.01756f
C650 CIN a_6741_2961# 0.00105f
C651 B a_1999_2695# 0.00187f
C652 a_13976_3192# a_14129_2675# -0
C653 a_16463_2943# COUT 0.00193f
C654 li_22548_2776# COUT 0
C655 a_14393_2675# A 0.00861f
C656 sky130_fd_sc_hs__inv_2_0/w_n38_332# COUT 0.00557f
C657 a_17568_3188# a_16463_2943# -0
C658 ua[1] VNB 0.1369f
C659 ua[2] VNB 0.1369f
C660 ua[3] VNB 0.1369f
C661 ua[4] VNB 0.1369f
C662 ua[5] VNB 0.1369f
C663 ua[6] VNB 0.1369f
C664 ua[7] VNB 0.1369f
C665 ena VNB 0.06503f
C666 clk VNB 0.03887f
C667 rst_n VNB 0.03887f
C668 ui_in[0] VNB 0.03887f
C669 ui_in[1] VNB 0.03887f
C670 ui_in[2] VNB 0.03887f
C671 ui_in[3] VNB 0.03887f
C672 ui_in[4] VNB 0.03887f
C673 ui_in[5] VNB 0.03887f
C674 ui_in[6] VNB 0.03887f
C675 ui_in[7] VNB 0.03887f
C676 uio_in[0] VNB 0.03887f
C677 uio_in[1] VNB 0.03887f
C678 uio_in[2] VNB 0.03887f
C679 uio_in[3] VNB 0.03887f
C680 uio_in[4] VNB 0.03887f
C681 uio_in[5] VNB 0.03887f
C682 uio_in[6] VNB 0.03887f
C683 uio_in[7] VNB 0.03887f
C684 uo_out[0] VNB 0.03887f
C685 uo_out[1] VNB 0.03887f
C686 uo_out[2] VNB 0.03887f
C687 uo_out[3] VNB 0.03887f
C688 uo_out[4] VNB 0.03887f
C689 uo_out[5] VNB 0.03887f
C690 uo_out[6] VNB 0.03887f
C691 uo_out[7] VNB 0.03887f
C692 uio_out[0] VNB 0.03887f
C693 uio_out[1] VNB 0.03887f
C694 uio_out[2] VNB 0.03887f
C695 uio_out[3] VNB 0.03887f
C696 uio_out[4] VNB 0.03887f
C697 uio_out[5] VNB 0.03887f
C698 uio_out[6] VNB 0.03887f
C699 uio_out[7] VNB 0.03887f
C700 uio_oe[0] VNB 0.03887f
C701 uio_oe[1] VNB 0.03887f
C702 uio_oe[2] VNB 0.03887f
C703 uio_oe[3] VNB 0.03887f
C704 uio_oe[4] VNB 0.03887f
C705 uio_oe[5] VNB 0.03887f
C706 uio_oe[6] VNB 0.03887f
C707 uio_oe[7] VNB 0.06503f
C708 a_17568_3188# VNB 0.30033f
C709 a_16038_3188# VNB 0.14774f
C710 a_15506_3192# VNB 0.2969f
C711 a_13976_3192# VNB 0.14781f
C712 a_13432_3194# VNB 0.29703f
C713 a_11902_3194# VNB 0.14774f
C714 a_11370_3198# VNB 0.27898f
C715 a_9840_3198# VNB 0.1477f
C716 a_9310_3202# VNB 0.29686f
C717 a_7780_3202# VNB 0.14774f
C718 a_7248_3206# VNB 0.2969f
C719 a_5718_3206# VNB 0.14781f
C720 B VNB 37.25793f
C721 a_5174_3208# VNB 0.29703f
C722 a_3644_3208# VNB 0.14774f
C723 a_3112_3212# VNB 0.2969f
C724 CIN VNB 2.22921f
C725 a_1582_3212# VNB 0.15472f
C726 COUT VNB 4.90409f
C727 a_17054_2671# VNB 0.01137f
C728 a_16455_2671# VNB 0.00504f
C729 a_17061_2943# VNB 0.00204f
C730 a_16463_2943# VNB 0.00129f
C731 ua[0] VNB 2.07042f
C732 w_28060_2795# VNB 1.49072f
C733 sky130_fd_sc_hs__fa_1_2/CIN VNB 0.50058f
C734 sky130_fd_sc_hs__fa_1_3/CIN VNB 0.50559f
C735 a_6734_2689# VNB 0.01137f
C736 a_6135_2689# VNB 0.00504f
C737 a_6741_2961# VNB 0.00204f
C738 a_6143_2961# VNB 0.00129f
C739 sky130_fd_sc_hs__fa_1_5/CIN VNB 0.40472f
C740 a_14992_2675# VNB 0.01137f
C741 a_14393_2675# VNB 0.00504f
C742 a_14999_2947# VNB 0.00204f
C743 a_14401_2947# VNB 0.00129f
C744 a_29450_3031# VNB 1.72277f
C745 w_26254_2813# VNB 1.49072f
C746 a_8796_2685# VNB 0.01137f
C747 a_8197_2685# VNB 0.00504f
C748 a_8803_2957# VNB 0.00204f
C749 a_8205_2957# VNB 0.00129f
C750 w_18084_2861# VNB 0.33898f
C751 sky130_fd_sc_hd__inv_1_0/w_n38_261# VNB 0.33898f
C752 a_27644_3049# VNB 1.71743f
C753 sky130_fd_sc_hd__inv_16_0/w_n38_261# VNB 1.49072f
C754 a_4660_2691# VNB 0.01137f
C755 a_4061_2691# VNB 0.00504f
C756 a_4667_2963# VNB 0.00204f
C757 a_4069_2963# VNB 0.00129f
C758 sky130_fd_sc_hs__inv_2_0/w_n38_332# VNB 0.40622f
C759 sky130_fd_sc_hs__fa_1_1/CIN VNB 0.50093f
C760 A VNB 40.0673f
C761 SUM VNB 0.61793f
C762 VPB VNB 16.70885f
C763 a_2598_2695# VNB 0.01137f
C764 a_1999_2695# VNB 0.00504f
C765 a_2605_2967# VNB 0.00204f
C766 a_2007_2967# VNB 0.00129f
C767 sky130_fd_sc_hd__inv_2_0/w_n38_261# VNB 0.33898f
C768 sky130_fd_sc_hd__inv_4_0/w_n38_261# VNB 0.51617f
C769 li_21382_2780# VNB 0.97225f
C770 sky130_fd_sc_hd__inv_6_0/w_n38_261# VNB 0.69336f
C771 li_24080_2768# VNB 1.76222f
C772 sky130_fd_sc_hd__inv_12_0/w_n38_261# VNB 1.22494f
C773 li_22548_2776# VNB 1.35117f
C774 sky130_fd_sc_hd__inv_8_0/w_n38_261# VNB 0.87055f
C775 sky130_fd_sc_hs__fa_1_6/CIN VNB 0.51989f
C776 sky130_fd_sc_hs__fa_1_7/CIN VNB 0.51916f
C777 a_10856_2681# VNB 0.01137f
C778 a_10257_2681# VNB 0.00504f
C779 a_10863_2953# VNB 0.00204f
C780 a_10265_2953# VNB 0.00129f
C781 sky130_fd_sc_hs__fa_1_4/CIN VNB 0.52445f
C782 a_12918_2677# VNB 0.01137f
C783 a_12319_2677# VNB 0.00504f
C784 a_12925_2949# VNB 0.00204f
C785 a_12327_2949# VNB 0.00129f
.ends

